module hardware_wrapper(
    
)