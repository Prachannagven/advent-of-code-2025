`timescale 1ns/1ps

module zero_counter_tb;

    // DUT inputs
    reg  [31:0] data_in;
    reg         dir_r;
    reg         clk;
    reg         rst;

    // DUT output
    wire [15:0] zero_count;
    wire [15:0] zero_cross;

    // Instantiate DUT
    zero_counter dut (
        .data_in(data_in),
        .dir_r(dir_r),
        .clk(clk),
        .rst(rst),
        .zero_count(zero_count),
        .zero_cross(zero_cross)
    );

    // Clock: 10ns period = 100MHz
    always #5 clk = ~clk;

    // MAIN TEST
    initial begin
        // VCD dump for waveforms
        $dumpfile("zero_counter.vcd");
        $dumpvars(0, zero_counter_tb);

        $display("=== ZERO COUNTER TESTBENCH START ===");

        // Initialize signals
        clk     = 0;
        rst     = 0;
        data_in = 0;
        dir_r   = 0;

        // Reset pulse
        rst = 1;
        #20;
        rst = 0;

        // === BEGIN INPUT SEQUENCE ===
        @(posedge clk); dir_r = 0; data_in = 5;
        @(posedge clk); dir_r = 0; data_in = 37;
        @(posedge clk); dir_r = 0; data_in = 32;
        @(posedge clk); dir_r = 1; data_in = 5;
        @(posedge clk); dir_r = 0; data_in = 36;
        @(posedge clk); dir_r = 0; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 13;
        @(posedge clk); dir_r = 1; data_in = 17;
        @(posedge clk); dir_r = 0; data_in = 19;
        @(posedge clk); dir_r = 0; data_in = 34;
        @(posedge clk); dir_r = 1; data_in = 2;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 1; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 1; data_in = 35;
        @(posedge clk); dir_r = 1; data_in = 26;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 19;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 1; data_in = 10;
        @(posedge clk); dir_r = 0; data_in = 14;
        @(posedge clk); dir_r = 1; data_in = 43;
        @(posedge clk); dir_r = 1; data_in = 35;
        @(posedge clk); dir_r = 0; data_in = 25;
        @(posedge clk); dir_r = 0; data_in = 35;
        @(posedge clk); dir_r = 0; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 34;
        @(posedge clk); dir_r = 0; data_in = 3;
        @(posedge clk); dir_r = 1; data_in = 25;
        @(posedge clk); dir_r = 1; data_in = 7;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 1; data_in = 22;
        @(posedge clk); dir_r = 0; data_in = 19;
        @(posedge clk); dir_r = 0; data_in = 39;
        @(posedge clk); dir_r = 0; data_in = 24;
        @(posedge clk); dir_r = 0; data_in = 50;
        @(posedge clk); dir_r = 1; data_in = 30;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 39;
        @(posedge clk); dir_r = 1; data_in = 30;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 46;
        @(posedge clk); dir_r = 1; data_in = 45;
        @(posedge clk); dir_r = 0; data_in = 32;
        @(posedge clk); dir_r = 1; data_in = 22;
        @(posedge clk); dir_r = 1; data_in = 35;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 32;
        @(posedge clk); dir_r = 1; data_in = 32;
        @(posedge clk); dir_r = 1; data_in = 86;
        @(posedge clk); dir_r = 0; data_in = 67;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 34;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 1; data_in = 66;
        @(posedge clk); dir_r = 1; data_in = 34;
        @(posedge clk); dir_r = 1; data_in = 38;
        @(posedge clk); dir_r = 1; data_in = 33;
        @(posedge clk); dir_r = 0; data_in = 71;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 1; data_in = 91;
        @(posedge clk); dir_r = 1; data_in = 19;
        @(posedge clk); dir_r = 1; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 64;
        @(posedge clk); dir_r = 1; data_in = 36;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 1; data_in = 2;
        @(posedge clk); dir_r = 0; data_in = 45;
        @(posedge clk); dir_r = 0; data_in = 68;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 0; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 0; data_in = 35;
        @(posedge clk); dir_r = 0; data_in = 96;
        @(posedge clk); dir_r = 1; data_in = 41;
        @(posedge clk); dir_r = 1; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 93;
        @(posedge clk); dir_r = 0; data_in = 93;
        @(posedge clk); dir_r = 0; data_in = 8;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 16;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 54;
        @(posedge clk); dir_r = 0; data_in = 10;
        @(posedge clk); dir_r = 1; data_in = 14;
        @(posedge clk); dir_r = 1; data_in = 41;
        @(posedge clk); dir_r = 1; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 62;
        @(posedge clk); dir_r = 1; data_in = 89;
        @(posedge clk); dir_r = 1; data_in = 77;
        @(posedge clk); dir_r = 1; data_in = 13;
        @(posedge clk); dir_r = 0; data_in = 55;
        @(posedge clk); dir_r = 0; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 56;
        @(posedge clk); dir_r = 0; data_in = 56;
        @(posedge clk); dir_r = 0; data_in = 28;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 0; data_in = 28;
        @(posedge clk); dir_r = 0; data_in = 40;
        @(posedge clk); dir_r = 1; data_in = 427;
        @(posedge clk); dir_r = 0; data_in = 340;
        @(posedge clk); dir_r = 0; data_in = 75;
        @(posedge clk); dir_r = 1; data_in = 82;
        @(posedge clk); dir_r = 0; data_in = 2;
        @(posedge clk); dir_r = 0; data_in = 80;
        @(posedge clk); dir_r = 1; data_in = 926;
        @(posedge clk); dir_r = 1; data_in = 74;
        @(posedge clk); dir_r = 0; data_in = 846;
        @(posedge clk); dir_r = 1; data_in = 29;
        @(posedge clk); dir_r = 0; data_in = 13;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 0; data_in = 15;
        @(posedge clk); dir_r = 0; data_in = 828;
        @(posedge clk); dir_r = 1; data_in = 75;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 0; data_in = 888;
        @(posedge clk); dir_r = 1; data_in = 25;
        @(posedge clk); dir_r = 0; data_in = 632;
        @(posedge clk); dir_r = 0; data_in = 86;
        @(posedge clk); dir_r = 0; data_in = 93;
        @(posedge clk); dir_r = 1; data_in = 51;
        @(posedge clk); dir_r = 0; data_in = 708;
        @(posedge clk); dir_r = 1; data_in = 409;
        @(posedge clk); dir_r = 1; data_in = 41;
        @(posedge clk); dir_r = 0; data_in = 55;
        @(posedge clk); dir_r = 0; data_in = 5;
        @(posedge clk); dir_r = 1; data_in = 460;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 0; data_in = 60;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 12;
        @(posedge clk); dir_r = 0; data_in = 230;
        @(posedge clk); dir_r = 1; data_in = 85;
        @(posedge clk); dir_r = 0; data_in = 3;
        @(posedge clk); dir_r = 0; data_in = 63;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 13;
        @(posedge clk); dir_r = 0; data_in = 80;
        @(posedge clk); dir_r = 0; data_in = 43;
        @(posedge clk); dir_r = 1; data_in = 23;
        @(posedge clk); dir_r = 0; data_in = 14;
        @(posedge clk); dir_r = 0; data_in = 86;
        @(posedge clk); dir_r = 1; data_in = 60;
        @(posedge clk); dir_r = 0; data_in = 60;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 82;
        @(posedge clk); dir_r = 1; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 26;
        @(posedge clk); dir_r = 0; data_in = 18;
        @(posedge clk); dir_r = 0; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 56;
        @(posedge clk); dir_r = 0; data_in = 96;
        @(posedge clk); dir_r = 0; data_in = 277;
        @(posedge clk); dir_r = 1; data_in = 77;
        @(posedge clk); dir_r = 1; data_in = 88;
        @(posedge clk); dir_r = 1; data_in = 212;
        @(posedge clk); dir_r = 1; data_in = 471;
        @(posedge clk); dir_r = 0; data_in = 77;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 96;
        @(posedge clk); dir_r = 1; data_in = 38;
        @(posedge clk); dir_r = 1; data_in = 66;
        @(posedge clk); dir_r = 1; data_in = 83;
        @(posedge clk); dir_r = 0; data_in = 29;
        @(posedge clk); dir_r = 0; data_in = 54;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 62;
        @(posedge clk); dir_r = 0; data_in = 6;
        @(posedge clk); dir_r = 0; data_in = 5;
        @(posedge clk); dir_r = 1; data_in = 401;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 0; data_in = 192;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 0; data_in = 615;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 0; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 33;
        @(posedge clk); dir_r = 1; data_in = 94;
        @(posedge clk); dir_r = 1; data_in = 50;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 94;
        @(posedge clk); dir_r = 0; data_in = 163;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 0; data_in = 91;
        @(posedge clk); dir_r = 1; data_in = 273;
        @(posedge clk); dir_r = 1; data_in = 83;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 3;
        @(posedge clk); dir_r = 1; data_in = 17;
        @(posedge clk); dir_r = 0; data_in = 85;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 1; data_in = 61;
        @(posedge clk); dir_r = 1; data_in = 63;
        @(posedge clk); dir_r = 1; data_in = 537;
        @(posedge clk); dir_r = 0; data_in = 395;
        @(posedge clk); dir_r = 0; data_in = 5;
        @(posedge clk); dir_r = 1; data_in = 297;
        @(posedge clk); dir_r = 0; data_in = 97;
        @(posedge clk); dir_r = 0; data_in = 194;
        @(posedge clk); dir_r = 0; data_in = 806;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 127;
        @(posedge clk); dir_r = 0; data_in = 879;
        @(posedge clk); dir_r = 0; data_in = 164;
        @(posedge clk); dir_r = 0; data_in = 56;
        @(posedge clk); dir_r = 0; data_in = 95;
        @(posedge clk); dir_r = 0; data_in = 62;
        @(posedge clk); dir_r = 0; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 183;
        @(posedge clk); dir_r = 0; data_in = 50;
        @(posedge clk); dir_r = 1; data_in = 25;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 0; data_in = 7;
        @(posedge clk); dir_r = 0; data_in = 80;
        @(posedge clk); dir_r = 1; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 6;
        @(posedge clk); dir_r = 0; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 74;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 40;
        @(posedge clk); dir_r = 1; data_in = 7;
        @(posedge clk); dir_r = 0; data_in = 67;
        @(posedge clk); dir_r = 1; data_in = 380;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 91;
        @(posedge clk); dir_r = 1; data_in = 83;
        @(posedge clk); dir_r = 0; data_in = 14;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 1; data_in = 10;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 1; data_in = 40;
        @(posedge clk); dir_r = 0; data_in = 40;
        @(posedge clk); dir_r = 0; data_in = 74;
        @(posedge clk); dir_r = 1; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 17;
        @(posedge clk); dir_r = 0; data_in = 74;
        @(posedge clk); dir_r = 0; data_in = 52;
        @(posedge clk); dir_r = 1; data_in = 96;
        @(posedge clk); dir_r = 0; data_in = 879;
        @(posedge clk); dir_r = 0; data_in = 7;
        @(posedge clk); dir_r = 0; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 173;
        @(posedge clk); dir_r = 0; data_in = 14;
        @(posedge clk); dir_r = 0; data_in = 66;
        @(posedge clk); dir_r = 1; data_in = 88;
        @(posedge clk); dir_r = 1; data_in = 25;
        @(posedge clk); dir_r = 1; data_in = 85;
        @(posedge clk); dir_r = 1; data_in = 867;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 1; data_in = 46;
        @(posedge clk); dir_r = 1; data_in = 30;
        @(posedge clk); dir_r = 1; data_in = 30;
        @(posedge clk); dir_r = 1; data_in = 486;
        @(posedge clk); dir_r = 0; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 150;
        @(posedge clk); dir_r = 1; data_in = 88;
        @(posedge clk); dir_r = 1; data_in = 85;
        @(posedge clk); dir_r = 1; data_in = 27;
        @(posedge clk); dir_r = 1; data_in = 726;
        @(posedge clk); dir_r = 0; data_in = 95;
        @(posedge clk); dir_r = 1; data_in = 55;
        @(posedge clk); dir_r = 0; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 7;
        @(posedge clk); dir_r = 0; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 32;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 1; data_in = 28;
        @(posedge clk); dir_r = 1; data_in = 599;
        @(posedge clk); dir_r = 1; data_in = 72;
        @(posedge clk); dir_r = 1; data_in = 37;
        @(posedge clk); dir_r = 1; data_in = 961;
        @(posedge clk); dir_r = 1; data_in = 30;
        @(posedge clk); dir_r = 1; data_in = 177;
        @(posedge clk); dir_r = 0; data_in = 8;
        @(posedge clk); dir_r = 0; data_in = 66;
        @(posedge clk); dir_r = 1; data_in = 99;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 1; data_in = 805;
        @(posedge clk); dir_r = 0; data_in = 52;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 64;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 37;
        @(posedge clk); dir_r = 0; data_in = 17;
        @(posedge clk); dir_r = 1; data_in = 520;
        @(posedge clk); dir_r = 0; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 1; data_in = 91;
        @(posedge clk); dir_r = 0; data_in = 69;
        @(posedge clk); dir_r = 0; data_in = 56;
        @(posedge clk); dir_r = 0; data_in = 55;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 54;
        @(posedge clk); dir_r = 0; data_in = 429;
        @(posedge clk); dir_r = 1; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 58;
        @(posedge clk); dir_r = 1; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 43;
        @(posedge clk); dir_r = 0; data_in = 504;
        @(posedge clk); dir_r = 0; data_in = 159;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 32;
        @(posedge clk); dir_r = 0; data_in = 17;
        @(posedge clk); dir_r = 1; data_in = 62;
        @(posedge clk); dir_r = 0; data_in = 46;
        @(posedge clk); dir_r = 0; data_in = 47;
        @(posedge clk); dir_r = 1; data_in = 392;
        @(posedge clk); dir_r = 1; data_in = 36;
        @(posedge clk); dir_r = 1; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 562;
        @(posedge clk); dir_r = 0; data_in = 22;
        @(posedge clk); dir_r = 0; data_in = 46;
        @(posedge clk); dir_r = 0; data_in = 8;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 22;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 1; data_in = 78;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 0; data_in = 86;
        @(posedge clk); dir_r = 0; data_in = 764;
        @(posedge clk); dir_r = 0; data_in = 97;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 1; data_in = 39;
        @(posedge clk); dir_r = 1; data_in = 982;
        @(posedge clk); dir_r = 0; data_in = 75;
        @(posedge clk); dir_r = 1; data_in = 240;
        @(posedge clk); dir_r = 1; data_in = 77;
        @(posedge clk); dir_r = 1; data_in = 57;
        @(posedge clk); dir_r = 1; data_in = 28;
        @(posedge clk); dir_r = 0; data_in = 86;
        @(posedge clk); dir_r = 0; data_in = 28;
        @(posedge clk); dir_r = 0; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 357;
        @(posedge clk); dir_r = 1; data_in = 64;
        @(posedge clk); dir_r = 1; data_in = 93;
        @(posedge clk); dir_r = 0; data_in = 462;
        @(posedge clk); dir_r = 0; data_in = 82;
        @(posedge clk); dir_r = 1; data_in = 93;
        @(posedge clk); dir_r = 1; data_in = 7;
        @(posedge clk); dir_r = 0; data_in = 6;
        @(posedge clk); dir_r = 0; data_in = 50;
        @(posedge clk); dir_r = 1; data_in = 77;
        @(posedge clk); dir_r = 0; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 60;
        @(posedge clk); dir_r = 1; data_in = 18;
        @(posedge clk); dir_r = 1; data_in = 60;
        @(posedge clk); dir_r = 0; data_in = 78;
        @(posedge clk); dir_r = 0; data_in = 545;
        @(posedge clk); dir_r = 1; data_in = 45;
        @(posedge clk); dir_r = 0; data_in = 303;
        @(posedge clk); dir_r = 0; data_in = 46;
        @(posedge clk); dir_r = 0; data_in = 51;
        @(posedge clk); dir_r = 1; data_in = 94;
        @(posedge clk); dir_r = 0; data_in = 8;
        @(posedge clk); dir_r = 1; data_in = 492;
        @(posedge clk); dir_r = 1; data_in = 48;
        @(posedge clk); dir_r = 1; data_in = 185;
        @(posedge clk); dir_r = 0; data_in = 51;
        @(posedge clk); dir_r = 0; data_in = 28;
        @(posedge clk); dir_r = 1; data_in = 14;
        @(posedge clk); dir_r = 0; data_in = 353;
        @(posedge clk); dir_r = 0; data_in = 25;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 0; data_in = 868;
        @(posedge clk); dir_r = 1; data_in = 982;
        @(posedge clk); dir_r = 0; data_in = 30;
        @(posedge clk); dir_r = 0; data_in = 82;
        @(posedge clk); dir_r = 0; data_in = 25;
        @(posedge clk); dir_r = 1; data_in = 543;
        @(posedge clk); dir_r = 0; data_in = 828;
        @(posedge clk); dir_r = 0; data_in = 60;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 0; data_in = 19;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 85;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 30;
        @(posedge clk); dir_r = 1; data_in = 855;
        @(posedge clk); dir_r = 0; data_in = 18;
        @(posedge clk); dir_r = 0; data_in = 82;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 112;
        @(posedge clk); dir_r = 0; data_in = 940;
        @(posedge clk); dir_r = 0; data_in = 31;
        @(posedge clk); dir_r = 1; data_in = 327;
        @(posedge clk); dir_r = 1; data_in = 48;
        @(posedge clk); dir_r = 0; data_in = 3;
        @(posedge clk); dir_r = 0; data_in = 75;
        @(posedge clk); dir_r = 1; data_in = 93;
        @(posedge clk); dir_r = 0; data_in = 2;
        @(posedge clk); dir_r = 0; data_in = 35;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 1; data_in = 198;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 1; data_in = 69;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 290;
        @(posedge clk); dir_r = 1; data_in = 64;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 72;
        @(posedge clk); dir_r = 1; data_in = 89;
        @(posedge clk); dir_r = 0; data_in = 54;
        @(posedge clk); dir_r = 0; data_in = 243;
        @(posedge clk); dir_r = 0; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 414;
        @(posedge clk); dir_r = 1; data_in = 23;
        @(posedge clk); dir_r = 1; data_in = 39;
        @(posedge clk); dir_r = 1; data_in = 61;
        @(posedge clk); dir_r = 1; data_in = 91;
        @(posedge clk); dir_r = 0; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 41;
        @(posedge clk); dir_r = 0; data_in = 77;
        @(posedge clk); dir_r = 1; data_in = 273;
        @(posedge clk); dir_r = 0; data_in = 32;
        @(posedge clk); dir_r = 1; data_in = 59;
        @(posedge clk); dir_r = 0; data_in = 579;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 1; data_in = 46;
        @(posedge clk); dir_r = 0; data_in = 7;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 1; data_in = 80;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 88;
        @(posedge clk); dir_r = 0; data_in = 65;
        @(posedge clk); dir_r = 1; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 88;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 0; data_in = 33;
        @(posedge clk); dir_r = 1; data_in = 19;
        @(posedge clk); dir_r = 0; data_in = 57;
        @(posedge clk); dir_r = 1; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 1; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 442;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 37;
        @(posedge clk); dir_r = 0; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 376;
        @(posedge clk); dir_r = 1; data_in = 23;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 96;
        @(posedge clk); dir_r = 1; data_in = 43;
        @(posedge clk); dir_r = 0; data_in = 41;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 0; data_in = 124;
        @(posedge clk); dir_r = 0; data_in = 872;
        @(posedge clk); dir_r = 0; data_in = 54;
        @(posedge clk); dir_r = 1; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 19;
        @(posedge clk); dir_r = 0; data_in = 95;
        @(posedge clk); dir_r = 0; data_in = 15;
        @(posedge clk); dir_r = 0; data_in = 90;
        @(posedge clk); dir_r = 1; data_in = 920;
        @(posedge clk); dir_r = 0; data_in = 62;
        @(posedge clk); dir_r = 1; data_in = 43;
        @(posedge clk); dir_r = 1; data_in = 99;
        @(posedge clk); dir_r = 1; data_in = 3;
        @(posedge clk); dir_r = 0; data_in = 944;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 0; data_in = 106;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 0; data_in = 91;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 0; data_in = 35;
        @(posedge clk); dir_r = 1; data_in = 33;
        @(posedge clk); dir_r = 1; data_in = 61;
        @(posedge clk); dir_r = 1; data_in = 52;
        @(posedge clk); dir_r = 0; data_in = 77;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 0; data_in = 33;
        @(posedge clk); dir_r = 1; data_in = 696;
        @(posedge clk); dir_r = 0; data_in = 19;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 77;
        @(posedge clk); dir_r = 0; data_in = 45;
        @(posedge clk); dir_r = 0; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 86;
        @(posedge clk); dir_r = 1; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 49;
        @(posedge clk); dir_r = 0; data_in = 1;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 35;
        @(posedge clk); dir_r = 0; data_in = 283;
        @(posedge clk); dir_r = 1; data_in = 48;
        @(posedge clk); dir_r = 0; data_in = 57;
        @(posedge clk); dir_r = 0; data_in = 38;
        @(posedge clk); dir_r = 1; data_in = 96;
        @(posedge clk); dir_r = 0; data_in = 7;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 1; data_in = 247;
        @(posedge clk); dir_r = 1; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 24;
        @(posedge clk); dir_r = 0; data_in = 3;
        @(posedge clk); dir_r = 1; data_in = 77;
        @(posedge clk); dir_r = 1; data_in = 93;
        @(posedge clk); dir_r = 0; data_in = 93;
        @(posedge clk); dir_r = 0; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 1; data_in = 80;
        @(posedge clk); dir_r = 0; data_in = 46;
        @(posedge clk); dir_r = 0; data_in = 49;
        @(posedge clk); dir_r = 1; data_in = 697;
        @(posedge clk); dir_r = 1; data_in = 52;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 1; data_in = 95;
        @(posedge clk); dir_r = 1; data_in = 877;
        @(posedge clk); dir_r = 1; data_in = 59;
        @(posedge clk); dir_r = 0; data_in = 17;
        @(posedge clk); dir_r = 1; data_in = 25;
        @(posedge clk); dir_r = 1; data_in = 7;
        @(posedge clk); dir_r = 0; data_in = 792;
        @(posedge clk); dir_r = 0; data_in = 707;
        @(posedge clk); dir_r = 0; data_in = 55;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 1; data_in = 571;
        @(posedge clk); dir_r = 1; data_in = 74;
        @(posedge clk); dir_r = 1; data_in = 74;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 0; data_in = 794;
        @(posedge clk); dir_r = 1; data_in = 23;
        @(posedge clk); dir_r = 0; data_in = 94;
        @(posedge clk); dir_r = 1; data_in = 26;
        @(posedge clk); dir_r = 0; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 856;
        @(posedge clk); dir_r = 0; data_in = 515;
        @(posedge clk); dir_r = 1; data_in = 71;
        @(posedge clk); dir_r = 1; data_in = 88;
        @(posedge clk); dir_r = 0; data_in = 5;
        @(posedge clk); dir_r = 0; data_in = 732;
        @(posedge clk); dir_r = 0; data_in = 63;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 0; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 684;
        @(posedge clk); dir_r = 0; data_in = 10;
        @(posedge clk); dir_r = 1; data_in = 55;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 24;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 0; data_in = 909;
        @(posedge clk); dir_r = 1; data_in = 32;
        @(posedge clk); dir_r = 1; data_in = 705;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 84;
        @(posedge clk); dir_r = 0; data_in = 77;
        @(posedge clk); dir_r = 1; data_in = 48;
        @(posedge clk); dir_r = 1; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 56;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 0; data_in = 852;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 99;
        @(posedge clk); dir_r = 1; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 5;
        @(posedge clk); dir_r = 1; data_in = 258;
        @(posedge clk); dir_r = 0; data_in = 32;
        @(posedge clk); dir_r = 1; data_in = 32;
        @(posedge clk); dir_r = 0; data_in = 5;
        @(posedge clk); dir_r = 1; data_in = 46;
        @(posedge clk); dir_r = 0; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 446;
        @(posedge clk); dir_r = 0; data_in = 85;
        @(posedge clk); dir_r = 0; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 32;
        @(posedge clk); dir_r = 0; data_in = 51;
        @(posedge clk); dir_r = 1; data_in = 61;
        @(posedge clk); dir_r = 1; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 37;
        @(posedge clk); dir_r = 0; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 460;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 0; data_in = 39;
        @(posedge clk); dir_r = 1; data_in = 36;
        @(posedge clk); dir_r = 0; data_in = 93;
        @(posedge clk); dir_r = 0; data_in = 282;
        @(posedge clk); dir_r = 0; data_in = 95;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 26;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 23;
        @(posedge clk); dir_r = 1; data_in = 77;
        @(posedge clk); dir_r = 1; data_in = 71;
        @(posedge clk); dir_r = 1; data_in = 17;
        @(posedge clk); dir_r = 1; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 54;
        @(posedge clk); dir_r = 0; data_in = 70;
        @(posedge clk); dir_r = 0; data_in = 36;
        @(posedge clk); dir_r = 0; data_in = 41;
        @(posedge clk); dir_r = 1; data_in = 48;
        @(posedge clk); dir_r = 1; data_in = 752;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 67;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 333;
        @(posedge clk); dir_r = 0; data_in = 58;
        @(posedge clk); dir_r = 1; data_in = 28;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 0; data_in = 91;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 806;
        @(posedge clk); dir_r = 1; data_in = 77;
        @(posedge clk); dir_r = 1; data_in = 59;
        @(posedge clk); dir_r = 0; data_in = 93;
        @(posedge clk); dir_r = 0; data_in = 35;
        @(posedge clk); dir_r = 0; data_in = 813;
        @(posedge clk); dir_r = 1; data_in = 905;
        @(posedge clk); dir_r = 1; data_in = 25;
        @(posedge clk); dir_r = 1; data_in = 75;
        @(posedge clk); dir_r = 1; data_in = 48;
        @(posedge clk); dir_r = 1; data_in = 722;
        @(posedge clk); dir_r = 0; data_in = 50;
        @(posedge clk); dir_r = 0; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 99;
        @(posedge clk); dir_r = 1; data_in = 50;
        @(posedge clk); dir_r = 0; data_in = 16;
        @(posedge clk); dir_r = 0; data_in = 19;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 1; data_in = 7;
        @(posedge clk); dir_r = 0; data_in = 48;
        @(posedge clk); dir_r = 1; data_in = 62;
        @(posedge clk); dir_r = 1; data_in = 19;
        @(posedge clk); dir_r = 0; data_in = 65;
        @(posedge clk); dir_r = 1; data_in = 88;
        @(posedge clk); dir_r = 0; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 783;
        @(posedge clk); dir_r = 1; data_in = 62;
        @(posedge clk); dir_r = 1; data_in = 5;
        @(posedge clk); dir_r = 0; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 74;
        @(posedge clk); dir_r = 0; data_in = 50;
        @(posedge clk); dir_r = 0; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 630;
        @(posedge clk); dir_r = 0; data_in = 78;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 90;
        @(posedge clk); dir_r = 0; data_in = 11;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 0; data_in = 449;
        @(posedge clk); dir_r = 0; data_in = 51;
        @(posedge clk); dir_r = 1; data_in = 811;
        @(posedge clk); dir_r = 1; data_in = 89;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 64;
        @(posedge clk); dir_r = 0; data_in = 5;
        @(posedge clk); dir_r = 0; data_in = 26;
        @(posedge clk); dir_r = 1; data_in = 8;
        @(posedge clk); dir_r = 0; data_in = 62;
        @(posedge clk); dir_r = 0; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 567;
        @(posedge clk); dir_r = 1; data_in = 71;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 1; data_in = 22;
        @(posedge clk); dir_r = 0; data_in = 35;
        @(posedge clk); dir_r = 1; data_in = 804;
        @(posedge clk); dir_r = 1; data_in = 59;
        @(posedge clk); dir_r = 0; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 33;
        @(posedge clk); dir_r = 0; data_in = 97;
        @(posedge clk); dir_r = 0; data_in = 25;
        @(posedge clk); dir_r = 1; data_in = 781;
        @(posedge clk); dir_r = 0; data_in = 678;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 5;
        @(posedge clk); dir_r = 0; data_in = 552;
        @(posedge clk); dir_r = 0; data_in = 48;
        @(posedge clk); dir_r = 0; data_in = 30;
        @(posedge clk); dir_r = 0; data_in = 49;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 1; data_in = 96;
        @(posedge clk); dir_r = 1; data_in = 29;
        @(posedge clk); dir_r = 0; data_in = 2;
        @(posedge clk); dir_r = 1; data_in = 37;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 0; data_in = 767;
        @(posedge clk); dir_r = 1; data_in = 172;
        @(posedge clk); dir_r = 1; data_in = 852;
        @(posedge clk); dir_r = 1; data_in = 958;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 54;
        @(posedge clk); dir_r = 0; data_in = 13;
        @(posedge clk); dir_r = 0; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 95;
        @(posedge clk); dir_r = 1; data_in = 393;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 758;
        @(posedge clk); dir_r = 1; data_in = 64;
        @(posedge clk); dir_r = 1; data_in = 36;
        @(posedge clk); dir_r = 0; data_in = 76;
        @(posedge clk); dir_r = 1; data_in = 76;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 1; data_in = 86;
        @(posedge clk); dir_r = 0; data_in = 426;
        @(posedge clk); dir_r = 1; data_in = 93;
        @(posedge clk); dir_r = 0; data_in = 165;
        @(posedge clk); dir_r = 0; data_in = 82;
        @(posedge clk); dir_r = 0; data_in = 18;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 0; data_in = 65;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 0; data_in = 49;
        @(posedge clk); dir_r = 0; data_in = 45;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 62;
        @(posedge clk); dir_r = 1; data_in = 22;
        @(posedge clk); dir_r = 1; data_in = 89;
        @(posedge clk); dir_r = 1; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 91;
        @(posedge clk); dir_r = 1; data_in = 33;
        @(posedge clk); dir_r = 0; data_in = 46;
        @(posedge clk); dir_r = 0; data_in = 49;
        @(posedge clk); dir_r = 1; data_in = 62;
        @(posedge clk); dir_r = 0; data_in = 362;
        @(posedge clk); dir_r = 0; data_in = 57;
        @(posedge clk); dir_r = 0; data_in = 81;
        @(posedge clk); dir_r = 0; data_in = 914;
        @(posedge clk); dir_r = 0; data_in = 86;
        @(posedge clk); dir_r = 0; data_in = 57;
        @(posedge clk); dir_r = 1; data_in = 89;
        @(posedge clk); dir_r = 1; data_in = 668;
        @(posedge clk); dir_r = 0; data_in = 36;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 1; data_in = 8;
        @(posedge clk); dir_r = 0; data_in = 97;
        @(posedge clk); dir_r = 1; data_in = 53;
        @(posedge clk); dir_r = 1; data_in = 53;
        @(posedge clk); dir_r = 1; data_in = 76;
        @(posedge clk); dir_r = 0; data_in = 93;
        @(posedge clk); dir_r = 1; data_in = 23;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 1; data_in = 460;
        @(posedge clk); dir_r = 0; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 33;
        @(posedge clk); dir_r = 0; data_in = 47;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 0; data_in = 54;
        @(posedge clk); dir_r = 0; data_in = 66;
        @(posedge clk); dir_r = 0; data_in = 48;
        @(posedge clk); dir_r = 1; data_in = 52;
        @(posedge clk); dir_r = 0; data_in = 12;
        @(posedge clk); dir_r = 0; data_in = 56;
        @(posedge clk); dir_r = 1; data_in = 941;
        @(posedge clk); dir_r = 1; data_in = 76;
        @(posedge clk); dir_r = 1; data_in = 3;
        @(posedge clk); dir_r = 1; data_in = 884;
        @(posedge clk); dir_r = 0; data_in = 71;
        @(posedge clk); dir_r = 1; data_in = 772;
        @(posedge clk); dir_r = 1; data_in = 28;
        @(posedge clk); dir_r = 0; data_in = 780;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 26;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 0; data_in = 1;
        @(posedge clk); dir_r = 0; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 242;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 82;
        @(posedge clk); dir_r = 0; data_in = 82;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 1; data_in = 94;
        @(posedge clk); dir_r = 1; data_in = 509;
        @(posedge clk); dir_r = 1; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 3;
        @(posedge clk); dir_r = 1; data_in = 72;
        @(posedge clk); dir_r = 1; data_in = 69;
        @(posedge clk); dir_r = 0; data_in = 37;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 385;
        @(posedge clk); dir_r = 1; data_in = 208;
        @(posedge clk); dir_r = 1; data_in = 629;
        @(posedge clk); dir_r = 1; data_in = 88;
        @(posedge clk); dir_r = 0; data_in = 752;
        @(posedge clk); dir_r = 0; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 0; data_in = 4;
        @(posedge clk); dir_r = 0; data_in = 97;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 36;
        @(posedge clk); dir_r = 0; data_in = 865;
        @(posedge clk); dir_r = 1; data_in = 225;
        @(posedge clk); dir_r = 0; data_in = 904;
        @(posedge clk); dir_r = 1; data_in = 26;
        @(posedge clk); dir_r = 0; data_in = 38;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 1; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 33;
        @(posedge clk); dir_r = 1; data_in = 673;
        @(posedge clk); dir_r = 1; data_in = 507;
        @(posedge clk); dir_r = 0; data_in = 2;
        @(posedge clk); dir_r = 1; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 25;
        @(posedge clk); dir_r = 0; data_in = 35;
        @(posedge clk); dir_r = 1; data_in = 3;
        @(posedge clk); dir_r = 0; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 0; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 54;
        @(posedge clk); dir_r = 0; data_in = 29;
        @(posedge clk); dir_r = 0; data_in = 17;
        @(posedge clk); dir_r = 1; data_in = 61;
        @(posedge clk); dir_r = 0; data_in = 248;
        @(posedge clk); dir_r = 0; data_in = 8;
        @(posedge clk); dir_r = 1; data_in = 82;
        @(posedge clk); dir_r = 1; data_in = 231;
        @(posedge clk); dir_r = 1; data_in = 75;
        @(posedge clk); dir_r = 1; data_in = 3;
        @(posedge clk); dir_r = 1; data_in = 968;
        @(posedge clk); dir_r = 0; data_in = 64;
        @(posedge clk); dir_r = 0; data_in = 46;
        @(posedge clk); dir_r = 1; data_in = 493;
        @(posedge clk); dir_r = 0; data_in = 47;
        @(posedge clk); dir_r = 1; data_in = 26;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 909;
        @(posedge clk); dir_r = 0; data_in = 942;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 83;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 1; data_in = 54;
        @(posedge clk); dir_r = 0; data_in = 93;
        @(posedge clk); dir_r = 1; data_in = 30;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 596;
        @(posedge clk); dir_r = 1; data_in = 67;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 0; data_in = 95;
        @(posedge clk); dir_r = 0; data_in = 76;
        @(posedge clk); dir_r = 0; data_in = 29;
        @(posedge clk); dir_r = 0; data_in = 52;
        @(posedge clk); dir_r = 0; data_in = 32;
        @(posedge clk); dir_r = 0; data_in = 65;
        @(posedge clk); dir_r = 0; data_in = 15;
        @(posedge clk); dir_r = 0; data_in = 36;
        @(posedge clk); dir_r = 1; data_in = 18;
        @(posedge clk); dir_r = 1; data_in = 71;
        @(posedge clk); dir_r = 0; data_in = 56;
        @(posedge clk); dir_r = 1; data_in = 67;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 0; data_in = 88;
        @(posedge clk); dir_r = 1; data_in = 76;
        @(posedge clk); dir_r = 0; data_in = 75;
        @(posedge clk); dir_r = 1; data_in = 167;
        @(posedge clk); dir_r = 1; data_in = 2;
        @(posedge clk); dir_r = 0; data_in = 292;
        @(posedge clk); dir_r = 1; data_in = 99;
        @(posedge clk); dir_r = 0; data_in = 795;
        @(posedge clk); dir_r = 1; data_in = 99;
        @(posedge clk); dir_r = 1; data_in = 202;
        @(posedge clk); dir_r = 1; data_in = 88;
        @(posedge clk); dir_r = 1; data_in = 10;
        @(posedge clk); dir_r = 0; data_in = 99;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 739;
        @(posedge clk); dir_r = 0; data_in = 65;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 0; data_in = 318;
        @(posedge clk); dir_r = 1; data_in = 26;
        @(posedge clk); dir_r = 0; data_in = 63;
        @(posedge clk); dir_r = 1; data_in = 18;
        @(posedge clk); dir_r = 1; data_in = 41;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 30;
        @(posedge clk); dir_r = 0; data_in = 30;
        @(posedge clk); dir_r = 1; data_in = 33;
        @(posedge clk); dir_r = 0; data_in = 70;
        @(posedge clk); dir_r = 0; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 43;
        @(posedge clk); dir_r = 0; data_in = 345;
        @(posedge clk); dir_r = 1; data_in = 210;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 0; data_in = 374;
        @(posedge clk); dir_r = 0; data_in = 968;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 970;
        @(posedge clk); dir_r = 1; data_in = 436;
        @(posedge clk); dir_r = 0; data_in = 37;
        @(posedge clk); dir_r = 0; data_in = 99;
        @(posedge clk); dir_r = 0; data_in = 29;
        @(posedge clk); dir_r = 0; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 71;
        @(posedge clk); dir_r = 1; data_in = 571;
        @(posedge clk); dir_r = 1; data_in = 92;
        @(posedge clk); dir_r = 1; data_in = 40;
        @(posedge clk); dir_r = 0; data_in = 309;
        @(posedge clk); dir_r = 1; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 85;
        @(posedge clk); dir_r = 1; data_in = 67;
        @(posedge clk); dir_r = 0; data_in = 170;
        @(posedge clk); dir_r = 1; data_in = 35;
        @(posedge clk); dir_r = 1; data_in = 52;
        @(posedge clk); dir_r = 0; data_in = 69;
        @(posedge clk); dir_r = 0; data_in = 16;
        @(posedge clk); dir_r = 0; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 276;
        @(posedge clk); dir_r = 1; data_in = 89;
        @(posedge clk); dir_r = 0; data_in = 104;
        @(posedge clk); dir_r = 1; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 49;
        @(posedge clk); dir_r = 1; data_in = 949;
        @(posedge clk); dir_r = 1; data_in = 2;
        @(posedge clk); dir_r = 0; data_in = 861;
        @(posedge clk); dir_r = 0; data_in = 39;
        @(posedge clk); dir_r = 1; data_in = 67;
        @(posedge clk); dir_r = 0; data_in = 503;
        @(posedge clk); dir_r = 0; data_in = 564;
        @(posedge clk); dir_r = 0; data_in = 712;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 0; data_in = 84;
        @(posedge clk); dir_r = 0; data_in = 543;
        @(posedge clk); dir_r = 1; data_in = 80;
        @(posedge clk); dir_r = 0; data_in = 80;
        @(posedge clk); dir_r = 0; data_in = 25;
        @(posedge clk); dir_r = 0; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 269;
        @(posedge clk); dir_r = 0; data_in = 207;
        @(posedge clk); dir_r = 0; data_in = 78;
        @(posedge clk); dir_r = 0; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 358;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 0; data_in = 34;
        @(posedge clk); dir_r = 0; data_in = 85;
        @(posedge clk); dir_r = 1; data_in = 252;
        @(posedge clk); dir_r = 1; data_in = 75;
        @(posedge clk); dir_r = 1; data_in = 725;
        @(posedge clk); dir_r = 1; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 73;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 0; data_in = 57;
        @(posedge clk); dir_r = 1; data_in = 34;
        @(posedge clk); dir_r = 1; data_in = 43;
        @(posedge clk); dir_r = 0; data_in = 226;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 3;
        @(posedge clk); dir_r = 1; data_in = 775;
        @(posedge clk); dir_r = 0; data_in = 58;
        @(posedge clk); dir_r = 1; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 154;
        @(posedge clk); dir_r = 1; data_in = 46;
        @(posedge clk); dir_r = 0; data_in = 896;
        @(posedge clk); dir_r = 0; data_in = 72;
        @(posedge clk); dir_r = 1; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 46;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 940;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 837;
        @(posedge clk); dir_r = 1; data_in = 71;
        @(posedge clk); dir_r = 1; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 72;
        @(posedge clk); dir_r = 1; data_in = 98;
        @(posedge clk); dir_r = 1; data_in = 41;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 1; data_in = 865;
        @(posedge clk); dir_r = 1; data_in = 35;
        @(posedge clk); dir_r = 1; data_in = 173;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 1; data_in = 256;
        @(posedge clk); dir_r = 0; data_in = 37;
        @(posedge clk); dir_r = 1; data_in = 734;
        @(posedge clk); dir_r = 1; data_in = 58;
        @(posedge clk); dir_r = 1; data_in = 121;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 0; data_in = 22;
        @(posedge clk); dir_r = 0; data_in = 19;
        @(posedge clk); dir_r = 0; data_in = 19;
        @(posedge clk); dir_r = 0; data_in = 322;
        @(posedge clk); dir_r = 1; data_in = 13;
        @(posedge clk); dir_r = 0; data_in = 613;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 0; data_in = 34;
        @(posedge clk); dir_r = 1; data_in = 40;
        @(posedge clk); dir_r = 0; data_in = 40;
        @(posedge clk); dir_r = 0; data_in = 52;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 399;
        @(posedge clk); dir_r = 0; data_in = 57;
        @(posedge clk); dir_r = 1; data_in = 17;
        @(posedge clk); dir_r = 0; data_in = 156;
        @(posedge clk); dir_r = 1; data_in = 10;
        @(posedge clk); dir_r = 0; data_in = 32;
        @(posedge clk); dir_r = 1; data_in = 61;
        @(posedge clk); dir_r = 0; data_in = 97;
        @(posedge clk); dir_r = 0; data_in = 3;
        @(posedge clk); dir_r = 0; data_in = 380;
        @(posedge clk); dir_r = 0; data_in = 74;
        @(posedge clk); dir_r = 0; data_in = 19;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 30;
        @(posedge clk); dir_r = 1; data_in = 92;
        @(posedge clk); dir_r = 1; data_in = 334;
        @(posedge clk); dir_r = 0; data_in = 33;
        @(posedge clk); dir_r = 0; data_in = 93;
        @(posedge clk); dir_r = 0; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 7;
        @(posedge clk); dir_r = 0; data_in = 78;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 35;
        @(posedge clk); dir_r = 0; data_in = 937;
        @(posedge clk); dir_r = 0; data_in = 702;
        @(posedge clk); dir_r = 1; data_in = 3;
        @(posedge clk); dir_r = 0; data_in = 551;
        @(posedge clk); dir_r = 1; data_in = 61;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 34;
        @(posedge clk); dir_r = 0; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 94;
        @(posedge clk); dir_r = 0; data_in = 3;
        @(posedge clk); dir_r = 1; data_in = 43;
        @(posedge clk); dir_r = 0; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 54;
        @(posedge clk); dir_r = 1; data_in = 2;
        @(posedge clk); dir_r = 0; data_in = 35;
        @(posedge clk); dir_r = 1; data_in = 149;
        @(posedge clk); dir_r = 1; data_in = 714;
        @(posedge clk); dir_r = 0; data_in = 33;
        @(posedge clk); dir_r = 0; data_in = 30;
        @(posedge clk); dir_r = 1; data_in = 60;
        @(posedge clk); dir_r = 0; data_in = 99;
        @(posedge clk); dir_r = 1; data_in = 39;
        @(posedge clk); dir_r = 0; data_in = 94;
        @(posedge clk); dir_r = 1; data_in = 52;
        @(posedge clk); dir_r = 0; data_in = 33;
        @(posedge clk); dir_r = 1; data_in = 17;
        @(posedge clk); dir_r = 0; data_in = 268;
        @(posedge clk); dir_r = 1; data_in = 26;
        @(posedge clk); dir_r = 1; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 51;
        @(posedge clk); dir_r = 0; data_in = 757;
        @(posedge clk); dir_r = 0; data_in = 67;
        @(posedge clk); dir_r = 1; data_in = 95;
        @(posedge clk); dir_r = 0; data_in = 58;
        @(posedge clk); dir_r = 1; data_in = 99;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 312;
        @(posedge clk); dir_r = 1; data_in = 91;
        @(posedge clk); dir_r = 0; data_in = 67;
        @(posedge clk); dir_r = 0; data_in = 7;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 0; data_in = 85;
        @(posedge clk); dir_r = 0; data_in = 433;
        @(posedge clk); dir_r = 1; data_in = 618;
        @(posedge clk); dir_r = 0; data_in = 13;
        @(posedge clk); dir_r = 0; data_in = 66;
        @(posedge clk); dir_r = 0; data_in = 669;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 0; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 67;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 0; data_in = 68;
        @(posedge clk); dir_r = 0; data_in = 10;
        @(posedge clk); dir_r = 1; data_in = 878;
        @(posedge clk); dir_r = 1; data_in = 5;
        @(posedge clk); dir_r = 1; data_in = 64;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 973;
        @(posedge clk); dir_r = 0; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 56;
        @(posedge clk); dir_r = 1; data_in = 18;
        @(posedge clk); dir_r = 1; data_in = 773;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 0; data_in = 16;
        @(posedge clk); dir_r = 1; data_in = 2;
        @(posedge clk); dir_r = 0; data_in = 72;
        @(posedge clk); dir_r = 1; data_in = 46;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 1; data_in = 83;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 742;
        @(posedge clk); dir_r = 0; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 469;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 1; data_in = 13;
        @(posedge clk); dir_r = 0; data_in = 560;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 32;
        @(posedge clk); dir_r = 1; data_in = 41;
        @(posedge clk); dir_r = 1; data_in = 91;
        @(posedge clk); dir_r = 0; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 0; data_in = 43;
        @(posedge clk); dir_r = 1; data_in = 92;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 0; data_in = 19;
        @(posedge clk); dir_r = 1; data_in = 41;
        @(posedge clk); dir_r = 0; data_in = 538;
        @(posedge clk); dir_r = 1; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 38;
        @(posedge clk); dir_r = 0; data_in = 52;
        @(posedge clk); dir_r = 0; data_in = 10;
        @(posedge clk); dir_r = 0; data_in = 290;
        @(posedge clk); dir_r = 0; data_in = 34;
        @(posedge clk); dir_r = 0; data_in = 76;
        @(posedge clk); dir_r = 0; data_in = 40;
        @(posedge clk); dir_r = 0; data_in = 76;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 1; data_in = 95;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 62;
        @(posedge clk); dir_r = 1; data_in = 63;
        @(posedge clk); dir_r = 1; data_in = 51;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 509;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 0; data_in = 795;
        @(posedge clk); dir_r = 0; data_in = 719;
        @(posedge clk); dir_r = 0; data_in = 89;
        @(posedge clk); dir_r = 0; data_in = 19;
        @(posedge clk); dir_r = 1; data_in = 22;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 0; data_in = 14;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 1; data_in = 72;
        @(posedge clk); dir_r = 0; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 1; data_in = 50;
        @(posedge clk); dir_r = 1; data_in = 550;
        @(posedge clk); dir_r = 1; data_in = 769;
        @(posedge clk); dir_r = 0; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 657;
        @(posedge clk); dir_r = 1; data_in = 22;
        @(posedge clk); dir_r = 0; data_in = 50;
        @(posedge clk); dir_r = 0; data_in = 329;
        @(posedge clk); dir_r = 1; data_in = 664;
        @(posedge clk); dir_r = 1; data_in = 358;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 1; data_in = 4;
        @(posedge clk); dir_r = 0; data_in = 16;
        @(posedge clk); dir_r = 0; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 0; data_in = 66;
        @(posedge clk); dir_r = 1; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 679;
        @(posedge clk); dir_r = 1; data_in = 77;
        @(posedge clk); dir_r = 1; data_in = 22;
        @(posedge clk); dir_r = 0; data_in = 95;
        @(posedge clk); dir_r = 1; data_in = 95;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 0; data_in = 798;
        @(posedge clk); dir_r = 0; data_in = 36;
        @(posedge clk); dir_r = 1; data_in = 35;
        @(posedge clk); dir_r = 0; data_in = 74;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 1; data_in = 18;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 0; data_in = 62;
        @(posedge clk); dir_r = 0; data_in = 38;
        @(posedge clk); dir_r = 0; data_in = 30;
        @(posedge clk); dir_r = 0; data_in = 89;
        @(posedge clk); dir_r = 1; data_in = 19;
        @(posedge clk); dir_r = 1; data_in = 68;
        @(posedge clk); dir_r = 0; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 35;
        @(posedge clk); dir_r = 1; data_in = 50;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 0; data_in = 14;
        @(posedge clk); dir_r = 1; data_in = 78;
        @(posedge clk); dir_r = 0; data_in = 64;
        @(posedge clk); dir_r = 1; data_in = 58;
        @(posedge clk); dir_r = 0; data_in = 72;
        @(posedge clk); dir_r = 0; data_in = 86;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 4;
        @(posedge clk); dir_r = 0; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 57;
        @(posedge clk); dir_r = 0; data_in = 69;
        @(posedge clk); dir_r = 0; data_in = 267;
        @(posedge clk); dir_r = 0; data_in = 67;
        @(posedge clk); dir_r = 0; data_in = 33;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 0; data_in = 95;
        @(posedge clk); dir_r = 0; data_in = 66;
        @(posedge clk); dir_r = 1; data_in = 318;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 5;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 1; data_in = 2;
        @(posedge clk); dir_r = 1; data_in = 27;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 30;
        @(posedge clk); dir_r = 1; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 86;
        @(posedge clk); dir_r = 0; data_in = 153;
        @(posedge clk); dir_r = 1; data_in = 50;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 1; data_in = 86;
        @(posedge clk); dir_r = 1; data_in = 67;
        @(posedge clk); dir_r = 0; data_in = 85;
        @(posedge clk); dir_r = 1; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 71;
        @(posedge clk); dir_r = 1; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 18;
        @(posedge clk); dir_r = 0; data_in = 934;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 482;
        @(posedge clk); dir_r = 1; data_in = 328;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 979;
        @(posedge clk); dir_r = 1; data_in = 23;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 1; data_in = 28;
        @(posedge clk); dir_r = 0; data_in = 505;
        @(posedge clk); dir_r = 1; data_in = 23;
        @(posedge clk); dir_r = 1; data_in = 54;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 1; data_in = 57;
        @(posedge clk); dir_r = 0; data_in = 919;
        @(posedge clk); dir_r = 1; data_in = 60;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 1; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 27;
        @(posedge clk); dir_r = 0; data_in = 40;
        @(posedge clk); dir_r = 1; data_in = 36;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 0; data_in = 97;
        @(posedge clk); dir_r = 0; data_in = 898;
        @(posedge clk); dir_r = 0; data_in = 231;
        @(posedge clk); dir_r = 1; data_in = 798;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 948;
        @(posedge clk); dir_r = 1; data_in = 57;
        @(posedge clk); dir_r = 1; data_in = 389;
        @(posedge clk); dir_r = 0; data_in = 87;
        @(posedge clk); dir_r = 0; data_in = 834;
        @(posedge clk); dir_r = 0; data_in = 56;
        @(posedge clk); dir_r = 1; data_in = 845;
        @(posedge clk); dir_r = 1; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 1; data_in = 61;
        @(posedge clk); dir_r = 0; data_in = 561;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 1; data_in = 92;
        @(posedge clk); dir_r = 1; data_in = 7;
        @(posedge clk); dir_r = 0; data_in = 7;
        @(posedge clk); dir_r = 0; data_in = 2;
        @(posedge clk); dir_r = 1; data_in = 776;
        @(posedge clk); dir_r = 1; data_in = 526;
        @(posedge clk); dir_r = 1; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 1; data_in = 727;
        @(posedge clk); dir_r = 0; data_in = 60;
        @(posedge clk); dir_r = 0; data_in = 10;
        @(posedge clk); dir_r = 0; data_in = 50;
        @(posedge clk); dir_r = 0; data_in = 35;
        @(posedge clk); dir_r = 1; data_in = 735;
        @(posedge clk); dir_r = 0; data_in = 14;
        @(posedge clk); dir_r = 0; data_in = 686;
        @(posedge clk); dir_r = 0; data_in = 13;
        @(posedge clk); dir_r = 0; data_in = 55;
        @(posedge clk); dir_r = 0; data_in = 252;
        @(posedge clk); dir_r = 0; data_in = 422;
        @(posedge clk); dir_r = 0; data_in = 143;
        @(posedge clk); dir_r = 0; data_in = 50;
        @(posedge clk); dir_r = 1; data_in = 27;
        @(posedge clk); dir_r = 0; data_in = 398;
        @(posedge clk); dir_r = 0; data_in = 8;
        @(posedge clk); dir_r = 1; data_in = 443;
        @(posedge clk); dir_r = 1; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 0; data_in = 31;
        @(posedge clk); dir_r = 1; data_in = 63;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 632;
        @(posedge clk); dir_r = 1; data_in = 924;
        @(posedge clk); dir_r = 0; data_in = 32;
        @(posedge clk); dir_r = 1; data_in = 138;
        @(posedge clk); dir_r = 0; data_in = 70;
        @(posedge clk); dir_r = 0; data_in = 647;
        @(posedge clk); dir_r = 0; data_in = 55;
        @(posedge clk); dir_r = 0; data_in = 85;
        @(posedge clk); dir_r = 0; data_in = 85;
        @(posedge clk); dir_r = 1; data_in = 43;
        @(posedge clk); dir_r = 0; data_in = 28;
        @(posedge clk); dir_r = 0; data_in = 38;
        @(posedge clk); dir_r = 1; data_in = 93;
        @(posedge clk); dir_r = 0; data_in = 17;
        @(posedge clk); dir_r = 1; data_in = 40;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 1; data_in = 62;
        @(posedge clk); dir_r = 0; data_in = 82;
        @(posedge clk); dir_r = 0; data_in = 772;
        @(posedge clk); dir_r = 0; data_in = 8;
        @(posedge clk); dir_r = 0; data_in = 790;
        @(posedge clk); dir_r = 0; data_in = 10;
        @(posedge clk); dir_r = 1; data_in = 934;
        @(posedge clk); dir_r = 1; data_in = 29;
        @(posedge clk); dir_r = 0; data_in = 817;
        @(posedge clk); dir_r = 1; data_in = 517;
        @(posedge clk); dir_r = 0; data_in = 41;
        @(posedge clk); dir_r = 0; data_in = 822;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 1; data_in = 635;
        @(posedge clk); dir_r = 1; data_in = 41;
        @(posedge clk); dir_r = 1; data_in = 999;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 0; data_in = 78;
        @(posedge clk); dir_r = 1; data_in = 94;
        @(posedge clk); dir_r = 0; data_in = 26;
        @(posedge clk); dir_r = 1; data_in = 99;
        @(posedge clk); dir_r = 1; data_in = 8;
        @(posedge clk); dir_r = 0; data_in = 95;
        @(posedge clk); dir_r = 1; data_in = 94;
        @(posedge clk); dir_r = 0; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 308;
        @(posedge clk); dir_r = 0; data_in = 28;
        @(posedge clk); dir_r = 1; data_in = 567;
        @(posedge clk); dir_r = 1; data_in = 53;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 67;
        @(posedge clk); dir_r = 1; data_in = 23;
        @(posedge clk); dir_r = 0; data_in = 932;
        @(posedge clk); dir_r = 0; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 209;
        @(posedge clk); dir_r = 1; data_in = 51;
        @(posedge clk); dir_r = 0; data_in = 29;
        @(posedge clk); dir_r = 0; data_in = 3;
        @(posedge clk); dir_r = 1; data_in = 7;
        @(posedge clk); dir_r = 1; data_in = 592;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 39;
        @(posedge clk); dir_r = 1; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 71;
        @(posedge clk); dir_r = 0; data_in = 665;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 48;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 1; data_in = 49;
        @(posedge clk); dir_r = 1; data_in = 51;
        @(posedge clk); dir_r = 1; data_in = 69;
        @(posedge clk); dir_r = 0; data_in = 66;
        @(posedge clk); dir_r = 1; data_in = 27;
        @(posedge clk); dir_r = 0; data_in = 52;
        @(posedge clk); dir_r = 0; data_in = 78;
        @(posedge clk); dir_r = 0; data_in = 378;
        @(posedge clk); dir_r = 1; data_in = 690;
        @(posedge clk); dir_r = 0; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 1;
        @(posedge clk); dir_r = 0; data_in = 18;
        @(posedge clk); dir_r = 1; data_in = 7;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 93;
        @(posedge clk); dir_r = 0; data_in = 30;
        @(posedge clk); dir_r = 1; data_in = 923;
        @(posedge clk); dir_r = 0; data_in = 759;
        @(posedge clk); dir_r = 0; data_in = 419;
        @(posedge clk); dir_r = 1; data_in = 78;
        @(posedge clk); dir_r = 0; data_in = 15;
        @(posedge clk); dir_r = 0; data_in = 96;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 0; data_in = 583;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 426;
        @(posedge clk); dir_r = 1; data_in = 46;
        @(posedge clk); dir_r = 1; data_in = 121;
        @(posedge clk); dir_r = 0; data_in = 49;
        @(posedge clk); dir_r = 0; data_in = 72;
        @(posedge clk); dir_r = 1; data_in = 517;
        @(posedge clk); dir_r = 1; data_in = 661;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 0; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 29;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 26;
        @(posedge clk); dir_r = 1; data_in = 40;
        @(posedge clk); dir_r = 1; data_in = 88;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 772;
        @(posedge clk); dir_r = 1; data_in = 51;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 88;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 0; data_in = 91;
        @(posedge clk); dir_r = 1; data_in = 91;
        @(posedge clk); dir_r = 0; data_in = 38;
        @(posedge clk); dir_r = 0; data_in = 52;
        @(posedge clk); dir_r = 0; data_in = 10;
        @(posedge clk); dir_r = 1; data_in = 94;
        @(posedge clk); dir_r = 1; data_in = 480;
        @(posedge clk); dir_r = 0; data_in = 152;
        @(posedge clk); dir_r = 1; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 40;
        @(posedge clk); dir_r = 1; data_in = 851;
        @(posedge clk); dir_r = 0; data_in = 5;
        @(posedge clk); dir_r = 1; data_in = 954;
        @(posedge clk); dir_r = 1; data_in = 51;
        @(posedge clk); dir_r = 0; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 1; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 950;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 1; data_in = 606;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 1; data_in = 78;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 297;
        @(posedge clk); dir_r = 1; data_in = 72;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 0; data_in = 372;
        @(posedge clk); dir_r = 1; data_in = 112;
        @(posedge clk); dir_r = 1; data_in = 86;
        @(posedge clk); dir_r = 0; data_in = 726;
        @(posedge clk); dir_r = 0; data_in = 486;
        @(posedge clk); dir_r = 0; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 99;
        @(posedge clk); dir_r = 1; data_in = 35;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 1; data_in = 98;
        @(posedge clk); dir_r = 1; data_in = 602;
        @(posedge clk); dir_r = 1; data_in = 58;
        @(posedge clk); dir_r = 0; data_in = 31;
        @(posedge clk); dir_r = 1; data_in = 14;
        @(posedge clk); dir_r = 1; data_in = 859;
        @(posedge clk); dir_r = 1; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 43;
        @(posedge clk); dir_r = 0; data_in = 91;
        @(posedge clk); dir_r = 1; data_in = 71;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 4;
        @(posedge clk); dir_r = 0; data_in = 523;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 0; data_in = 12;
        @(posedge clk); dir_r = 1; data_in = 8;
        @(posedge clk); dir_r = 1; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 196;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 0; data_in = 569;
        @(posedge clk); dir_r = 1; data_in = 94;
        @(posedge clk); dir_r = 1; data_in = 30;
        @(posedge clk); dir_r = 0; data_in = 37;
        @(posedge clk); dir_r = 0; data_in = 80;
        @(posedge clk); dir_r = 0; data_in = 43;
        @(posedge clk); dir_r = 0; data_in = 48;
        @(posedge clk); dir_r = 1; data_in = 808;
        @(posedge clk); dir_r = 1; data_in = 64;
        @(posedge clk); dir_r = 1; data_in = 73;
        @(posedge clk); dir_r = 0; data_in = 37;
        @(posedge clk); dir_r = 0; data_in = 536;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 0; data_in = 62;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 0; data_in = 602;
        @(posedge clk); dir_r = 0; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 893;
        @(posedge clk); dir_r = 1; data_in = 17;
        @(posedge clk); dir_r = 1; data_in = 76;
        @(posedge clk); dir_r = 0; data_in = 10;
        @(posedge clk); dir_r = 0; data_in = 57;
        @(posedge clk); dir_r = 0; data_in = 86;
        @(posedge clk); dir_r = 0; data_in = 76;
        @(posedge clk); dir_r = 0; data_in = 28;
        @(posedge clk); dir_r = 1; data_in = 82;
        @(posedge clk); dir_r = 1; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 94;
        @(posedge clk); dir_r = 0; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 1; data_in = 338;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 95;
        @(posedge clk); dir_r = 1; data_in = 255;
        @(posedge clk); dir_r = 1; data_in = 40;
        @(posedge clk); dir_r = 1; data_in = 14;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 599;
        @(posedge clk); dir_r = 1; data_in = 40;
        @(posedge clk); dir_r = 1; data_in = 48;
        @(posedge clk); dir_r = 1; data_in = 93;
        @(posedge clk); dir_r = 1; data_in = 51;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 0; data_in = 86;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 91;
        @(posedge clk); dir_r = 0; data_in = 65;
        @(posedge clk); dir_r = 1; data_in = 74;
        @(posedge clk); dir_r = 1; data_in = 22;
        @(posedge clk); dir_r = 1; data_in = 85;
        @(posedge clk); dir_r = 0; data_in = 19;
        @(posedge clk); dir_r = 0; data_in = 798;
        @(posedge clk); dir_r = 1; data_in = 922;
        @(posedge clk); dir_r = 1; data_in = 57;
        @(posedge clk); dir_r = 0; data_in = 76;
        @(posedge clk); dir_r = 0; data_in = 72;
        @(posedge clk); dir_r = 0; data_in = 41;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 89;
        @(posedge clk); dir_r = 1; data_in = 60;
        @(posedge clk); dir_r = 0; data_in = 60;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 89;
        @(posedge clk); dir_r = 1; data_in = 95;
        @(posedge clk); dir_r = 0; data_in = 423;
        @(posedge clk); dir_r = 1; data_in = 339;
        @(posedge clk); dir_r = 0; data_in = 74;
        @(posedge clk); dir_r = 0; data_in = 148;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 0; data_in = 12;
        @(posedge clk); dir_r = 0; data_in = 18;
        @(posedge clk); dir_r = 0; data_in = 91;
        @(posedge clk); dir_r = 0; data_in = 894;
        @(posedge clk); dir_r = 1; data_in = 8;
        @(posedge clk); dir_r = 0; data_in = 49;
        @(posedge clk); dir_r = 1; data_in = 505;
        @(posedge clk); dir_r = 0; data_in = 561;
        @(posedge clk); dir_r = 1; data_in = 99;
        @(posedge clk); dir_r = 0; data_in = 99;
        @(posedge clk); dir_r = 0; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 790;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 980;
        @(posedge clk); dir_r = 0; data_in = 31;
        @(posedge clk); dir_r = 0; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 37;
        @(posedge clk); dir_r = 1; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 34;
        @(posedge clk); dir_r = 0; data_in = 80;
        @(posedge clk); dir_r = 1; data_in = 80;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 27;
        @(posedge clk); dir_r = 0; data_in = 22;
        @(posedge clk); dir_r = 0; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 64;
        @(posedge clk); dir_r = 1; data_in = 61;
        @(posedge clk); dir_r = 0; data_in = 25;
        @(posedge clk); dir_r = 0; data_in = 753;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 1; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 41;
        @(posedge clk); dir_r = 0; data_in = 933;
        @(posedge clk); dir_r = 0; data_in = 87;
        @(posedge clk); dir_r = 0; data_in = 24;
        @(posedge clk); dir_r = 0; data_in = 557;
        @(posedge clk); dir_r = 1; data_in = 74;
        @(posedge clk); dir_r = 1; data_in = 463;
        @(posedge clk); dir_r = 1; data_in = 259;
        @(posedge clk); dir_r = 0; data_in = 38;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 721;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 0; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 60;
        @(posedge clk); dir_r = 1; data_in = 64;
        @(posedge clk); dir_r = 1; data_in = 13;
        @(posedge clk); dir_r = 0; data_in = 929;
        @(posedge clk); dir_r = 1; data_in = 98;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 496;
        @(posedge clk); dir_r = 0; data_in = 2;
        @(posedge clk); dir_r = 0; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 4;
        @(posedge clk); dir_r = 0; data_in = 34;
        @(posedge clk); dir_r = 1; data_in = 146;
        @(posedge clk); dir_r = 1; data_in = 54;
        @(posedge clk); dir_r = 0; data_in = 958;
        @(posedge clk); dir_r = 0; data_in = 64;
        @(posedge clk); dir_r = 1; data_in = 220;
        @(posedge clk); dir_r = 1; data_in = 32;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 32;
        @(posedge clk); dir_r = 1; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 49;
        @(posedge clk); dir_r = 0; data_in = 366;
        @(posedge clk); dir_r = 0; data_in = 56;
        @(posedge clk); dir_r = 1; data_in = 87;
        @(posedge clk); dir_r = 0; data_in = 96;
        @(posedge clk); dir_r = 0; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 63;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 987;
        @(posedge clk); dir_r = 0; data_in = 48;
        @(posedge clk); dir_r = 0; data_in = 650;
        @(posedge clk); dir_r = 1; data_in = 50;
        @(posedge clk); dir_r = 0; data_in = 54;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 1; data_in = 23;
        @(posedge clk); dir_r = 0; data_in = 46;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 0; data_in = 517;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 0; data_in = 484;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 0; data_in = 74;
        @(posedge clk); dir_r = 0; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 473;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 0; data_in = 41;
        @(posedge clk); dir_r = 0; data_in = 97;
        @(posedge clk); dir_r = 0; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 177;
        @(posedge clk); dir_r = 0; data_in = 504;
        @(posedge clk); dir_r = 0; data_in = 64;
        @(posedge clk); dir_r = 0; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 0; data_in = 71;
        @(posedge clk); dir_r = 0; data_in = 25;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 28;
        @(posedge clk); dir_r = 1; data_in = 48;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 62;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 13;
        @(posedge clk); dir_r = 0; data_in = 13;
        @(posedge clk); dir_r = 1; data_in = 695;
        @(posedge clk); dir_r = 0; data_in = 25;
        @(posedge clk); dir_r = 1; data_in = 43;
        @(posedge clk); dir_r = 1; data_in = 23;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 1; data_in = 28;
        @(posedge clk); dir_r = 0; data_in = 228;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 98;
        @(posedge clk); dir_r = 1; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 25;
        @(posedge clk); dir_r = 1; data_in = 51;
        @(posedge clk); dir_r = 0; data_in = 826;
        @(posedge clk); dir_r = 0; data_in = 1;
        @(posedge clk); dir_r = 0; data_in = 87;
        @(posedge clk); dir_r = 0; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 498;
        @(posedge clk); dir_r = 0; data_in = 13;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 1; data_in = 1;
        @(posedge clk); dir_r = 0; data_in = 55;
        @(posedge clk); dir_r = 0; data_in = 38;
        @(posedge clk); dir_r = 0; data_in = 7;
        @(posedge clk); dir_r = 1; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 204;
        @(posedge clk); dir_r = 0; data_in = 998;
        @(posedge clk); dir_r = 1; data_in = 80;
        @(posedge clk); dir_r = 0; data_in = 309;
        @(posedge clk); dir_r = 0; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 85;
        @(posedge clk); dir_r = 0; data_in = 47;
        @(posedge clk); dir_r = 1; data_in = 171;
        @(posedge clk); dir_r = 0; data_in = 39;
        @(posedge clk); dir_r = 1; data_in = 64;
        @(posedge clk); dir_r = 1; data_in = 336;
        @(posedge clk); dir_r = 0; data_in = 263;
        @(posedge clk); dir_r = 0; data_in = 76;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 0; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 74;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 1;
        @(posedge clk); dir_r = 0; data_in = 22;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 640;
        @(posedge clk); dir_r = 1; data_in = 204;
        @(posedge clk); dir_r = 1; data_in = 94;
        @(posedge clk); dir_r = 1; data_in = 93;
        @(posedge clk); dir_r = 1; data_in = 580;
        @(posedge clk); dir_r = 1; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 71;
        @(posedge clk); dir_r = 1; data_in = 50;
        @(posedge clk); dir_r = 1; data_in = 52;
        @(posedge clk); dir_r = 0; data_in = 54;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 376;
        @(posedge clk); dir_r = 1; data_in = 83;
        @(posedge clk); dir_r = 0; data_in = 66;
        @(posedge clk); dir_r = 0; data_in = 39;
        @(posedge clk); dir_r = 0; data_in = 2;
        @(posedge clk); dir_r = 0; data_in = 284;
        @(posedge clk); dir_r = 0; data_in = 28;
        @(posedge clk); dir_r = 0; data_in = 34;
        @(posedge clk); dir_r = 1; data_in = 58;
        @(posedge clk); dir_r = 0; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 17;
        @(posedge clk); dir_r = 0; data_in = 167;
        @(posedge clk); dir_r = 0; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 82;
        @(posedge clk); dir_r = 0; data_in = 88;
        @(posedge clk); dir_r = 0; data_in = 62;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 253;
        @(posedge clk); dir_r = 0; data_in = 35;
        @(posedge clk); dir_r = 0; data_in = 12;
        @(posedge clk); dir_r = 1; data_in = 113;
        @(posedge clk); dir_r = 0; data_in = 66;
        @(posedge clk); dir_r = 1; data_in = 96;
        @(posedge clk); dir_r = 0; data_in = 43;
        @(posedge clk); dir_r = 0; data_in = 95;
        @(posedge clk); dir_r = 1; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 0; data_in = 69;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 37;
        @(posedge clk); dir_r = 1; data_in = 810;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 1; data_in = 174;
        @(posedge clk); dir_r = 1; data_in = 1;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 0; data_in = 89;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 0; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 60;
        @(posedge clk); dir_r = 1; data_in = 18;
        @(posedge clk); dir_r = 1; data_in = 380;
        @(posedge clk); dir_r = 1; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 1; data_in = 684;
        @(posedge clk); dir_r = 1; data_in = 74;
        @(posedge clk); dir_r = 1; data_in = 26;
        @(posedge clk); dir_r = 0; data_in = 260;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 291;
        @(posedge clk); dir_r = 1; data_in = 95;
        @(posedge clk); dir_r = 1; data_in = 56;
        @(posedge clk); dir_r = 0; data_in = 81;
        @(posedge clk); dir_r = 0; data_in = 17;
        @(posedge clk); dir_r = 1; data_in = 86;
        @(posedge clk); dir_r = 1; data_in = 60;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 99;
        @(posedge clk); dir_r = 1; data_in = 82;
        @(posedge clk); dir_r = 1; data_in = 14;
        @(posedge clk); dir_r = 1; data_in = 56;
        @(posedge clk); dir_r = 0; data_in = 71;
        @(posedge clk); dir_r = 0; data_in = 29;
        @(posedge clk); dir_r = 0; data_in = 57;
        @(posedge clk); dir_r = 1; data_in = 757;
        @(posedge clk); dir_r = 1; data_in = 253;
        @(posedge clk); dir_r = 1; data_in = 947;
        @(posedge clk); dir_r = 1; data_in = 88;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 1; data_in = 73;
        @(posedge clk); dir_r = 0; data_in = 46;
        @(posedge clk); dir_r = 1; data_in = 40;
        @(posedge clk); dir_r = 0; data_in = 767;
        @(posedge clk); dir_r = 0; data_in = 76;
        @(posedge clk); dir_r = 1; data_in = 87;
        @(posedge clk); dir_r = 0; data_in = 58;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 1; data_in = 25;
        @(posedge clk); dir_r = 0; data_in = 25;
        @(posedge clk); dir_r = 0; data_in = 638;
        @(posedge clk); dir_r = 1; data_in = 13;
        @(posedge clk); dir_r = 1; data_in = 525;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 710;
        @(posedge clk); dir_r = 1; data_in = 779;
        @(posedge clk); dir_r = 0; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 138;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 0; data_in = 52;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 1; data_in = 482;
        @(posedge clk); dir_r = 0; data_in = 756;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 0; data_in = 30;
        @(posedge clk); dir_r = 1; data_in = 519;
        @(posedge clk); dir_r = 0; data_in = 280;
        @(posedge clk); dir_r = 0; data_in = 43;
        @(posedge clk); dir_r = 0; data_in = 66;
        @(posedge clk); dir_r = 0; data_in = 57;
        @(posedge clk); dir_r = 1; data_in = 58;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 1; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 36;
        @(posedge clk); dir_r = 0; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 66;
        @(posedge clk); dir_r = 0; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 82;
        @(posedge clk); dir_r = 1; data_in = 85;
        @(posedge clk); dir_r = 0; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 644;
        @(posedge clk); dir_r = 1; data_in = 941;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 0; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 26;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 26;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 235;
        @(posedge clk); dir_r = 0; data_in = 65;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 58;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 0; data_in = 39;
        @(posedge clk); dir_r = 1; data_in = 95;
        @(posedge clk); dir_r = 1; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 75;
        @(posedge clk); dir_r = 1; data_in = 85;
        @(posedge clk); dir_r = 0; data_in = 85;
        @(posedge clk); dir_r = 1; data_in = 99;
        @(posedge clk); dir_r = 0; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 0; data_in = 95;
        @(posedge clk); dir_r = 1; data_in = 95;
        @(posedge clk); dir_r = 0; data_in = 19;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 1; data_in = 75;
        @(posedge clk); dir_r = 1; data_in = 56;
        @(posedge clk); dir_r = 0; data_in = 26;
        @(posedge clk); dir_r = 1; data_in = 71;
        @(posedge clk); dir_r = 0; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 1; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 76;
        @(posedge clk); dir_r = 0; data_in = 41;
        @(posedge clk); dir_r = 1; data_in = 58;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 88;
        @(posedge clk); dir_r = 0; data_in = 945;
        @(posedge clk); dir_r = 0; data_in = 43;
        @(posedge clk); dir_r = 0; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 29;
        @(posedge clk); dir_r = 0; data_in = 551;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 27;
        @(posedge clk); dir_r = 1; data_in = 81;
        @(posedge clk); dir_r = 0; data_in = 14;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 0; data_in = 66;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 0; data_in = 844;
        @(posedge clk); dir_r = 0; data_in = 49;
        @(posedge clk); dir_r = 1; data_in = 56;
        @(posedge clk); dir_r = 1; data_in = 344;
        @(posedge clk); dir_r = 1; data_in = 54;
        @(posedge clk); dir_r = 1; data_in = 62;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 91;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 99;
        @(posedge clk); dir_r = 0; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 26;
        @(posedge clk); dir_r = 1; data_in = 76;
        @(posedge clk); dir_r = 1; data_in = 50;
        @(posedge clk); dir_r = 1; data_in = 860;
        @(posedge clk); dir_r = 1; data_in = 94;
        @(posedge clk); dir_r = 1; data_in = 923;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 0; data_in = 88;
        @(posedge clk); dir_r = 1; data_in = 83;
        @(posedge clk); dir_r = 0; data_in = 95;
        @(posedge clk); dir_r = 0; data_in = 12;
        @(posedge clk); dir_r = 0; data_in = 311;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 0; data_in = 33;
        @(posedge clk); dir_r = 1; data_in = 18;
        @(posedge clk); dir_r = 0; data_in = 18;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 36;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 0; data_in = 34;
        @(posedge clk); dir_r = 1; data_in = 75;
        @(posedge clk); dir_r = 1; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 630;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 1; data_in = 3;
        @(posedge clk); dir_r = 1; data_in = 95;
        @(posedge clk); dir_r = 0; data_in = 88;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 52;
        @(posedge clk); dir_r = 0; data_in = 49;
        @(posedge clk); dir_r = 0; data_in = 75;
        @(posedge clk); dir_r = 1; data_in = 17;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 10;
        @(posedge clk); dir_r = 0; data_in = 31;
        @(posedge clk); dir_r = 1; data_in = 61;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 10;
        @(posedge clk); dir_r = 0; data_in = 28;
        @(posedge clk); dir_r = 0; data_in = 878;
        @(posedge clk); dir_r = 1; data_in = 77;
        @(posedge clk); dir_r = 0; data_in = 381;
        @(posedge clk); dir_r = 0; data_in = 43;
        @(posedge clk); dir_r = 1; data_in = 43;
        @(posedge clk); dir_r = 1; data_in = 103;
        @(posedge clk); dir_r = 1; data_in = 35;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 1; data_in = 51;
        @(posedge clk); dir_r = 1; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 86;
        @(posedge clk); dir_r = 1; data_in = 61;
        @(posedge clk); dir_r = 1; data_in = 183;
        @(posedge clk); dir_r = 0; data_in = 66;
        @(posedge clk); dir_r = 1; data_in = 58;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 1; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 19;
        @(posedge clk); dir_r = 0; data_in = 919;
        @(posedge clk); dir_r = 1; data_in = 63;
        @(posedge clk); dir_r = 1; data_in = 37;
        @(posedge clk); dir_r = 0; data_in = 176;
        @(posedge clk); dir_r = 1; data_in = 27;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 33;
        @(posedge clk); dir_r = 1; data_in = 76;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 0; data_in = 56;
        @(posedge clk); dir_r = 0; data_in = 221;
        @(posedge clk); dir_r = 1; data_in = 620;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 1; data_in = 80;
        @(posedge clk); dir_r = 0; data_in = 906;
        @(posedge clk); dir_r = 1; data_in = 61;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 0; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 2;
        @(posedge clk); dir_r = 0; data_in = 633;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 1; data_in = 35;
        @(posedge clk); dir_r = 0; data_in = 8;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 1; data_in = 5;
        @(posedge clk); dir_r = 1; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 50;
        @(posedge clk); dir_r = 0; data_in = 95;
        @(posedge clk); dir_r = 0; data_in = 43;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 28;
        @(posedge clk); dir_r = 1; data_in = 791;
        @(posedge clk); dir_r = 0; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 399;
        @(posedge clk); dir_r = 1; data_in = 188;
        @(posedge clk); dir_r = 1; data_in = 28;
        @(posedge clk); dir_r = 0; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 97;
        @(posedge clk); dir_r = 1; data_in = 483;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 77;
        @(posedge clk); dir_r = 0; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 29;
        @(posedge clk); dir_r = 0; data_in = 54;
        @(posedge clk); dir_r = 1; data_in = 855;
        @(posedge clk); dir_r = 1; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 18;
        @(posedge clk); dir_r = 1; data_in = 846;
        @(posedge clk); dir_r = 0; data_in = 5;
        @(posedge clk); dir_r = 0; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 43;
        @(posedge clk); dir_r = 0; data_in = 13;
        @(posedge clk); dir_r = 0; data_in = 76;
        @(posedge clk); dir_r = 1; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 35;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 0; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 8;
        @(posedge clk); dir_r = 0; data_in = 224;
        @(posedge clk); dir_r = 0; data_in = 43;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 0; data_in = 85;
        @(posedge clk); dir_r = 0; data_in = 40;
        @(posedge clk); dir_r = 1; data_in = 29;
        @(posedge clk); dir_r = 0; data_in = 48;
        @(posedge clk); dir_r = 1; data_in = 778;
        @(posedge clk); dir_r = 1; data_in = 522;
        @(posedge clk); dir_r = 0; data_in = 235;
        @(posedge clk); dir_r = 0; data_in = 18;
        @(posedge clk); dir_r = 1; data_in = 553;
        @(posedge clk); dir_r = 0; data_in = 77;
        @(posedge clk); dir_r = 1; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 19;
        @(posedge clk); dir_r = 1; data_in = 577;
        @(posedge clk); dir_r = 1; data_in = 683;
        @(posedge clk); dir_r = 1; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 16;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 451;
        @(posedge clk); dir_r = 0; data_in = 51;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 931;
        @(posedge clk); dir_r = 1; data_in = 87;
        @(posedge clk); dir_r = 0; data_in = 86;
        @(posedge clk); dir_r = 0; data_in = 339;
        @(posedge clk); dir_r = 0; data_in = 46;
        @(posedge clk); dir_r = 0; data_in = 1;
        @(posedge clk); dir_r = 0; data_in = 202;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 0; data_in = 949;
        @(posedge clk); dir_r = 0; data_in = 25;
        @(posedge clk); dir_r = 0; data_in = 41;
        @(posedge clk); dir_r = 0; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 738;
        @(posedge clk); dir_r = 0; data_in = 81;
        @(posedge clk); dir_r = 0; data_in = 457;
        @(posedge clk); dir_r = 0; data_in = 74;
        @(posedge clk); dir_r = 1; data_in = 671;
        @(posedge clk); dir_r = 1; data_in = 76;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 624;
        @(posedge clk); dir_r = 1; data_in = 25;
        @(posedge clk); dir_r = 0; data_in = 51;
        @(posedge clk); dir_r = 0; data_in = 290;
        @(posedge clk); dir_r = 1; data_in = 94;
        @(posedge clk); dir_r = 1; data_in = 34;
        @(posedge clk); dir_r = 1; data_in = 656;
        @(posedge clk); dir_r = 1; data_in = 908;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 1; data_in = 40;
        @(posedge clk); dir_r = 0; data_in = 26;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 95;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 12;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 22;
        @(posedge clk); dir_r = 1; data_in = 71;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 0; data_in = 91;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 0; data_in = 65;
        @(posedge clk); dir_r = 1; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 57;
        @(posedge clk); dir_r = 0; data_in = 635;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 1; data_in = 27;
        @(posedge clk); dir_r = 0; data_in = 953;
        @(posedge clk); dir_r = 0; data_in = 570;
        @(posedge clk); dir_r = 0; data_in = 77;
        @(posedge clk); dir_r = 0; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 36;
        @(posedge clk); dir_r = 0; data_in = 928;
        @(posedge clk); dir_r = 1; data_in = 33;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 1; data_in = 99;
        @(posedge clk); dir_r = 0; data_in = 11;
        @(posedge clk); dir_r = 1; data_in = 26;
        @(posedge clk); dir_r = 1; data_in = 74;
        @(posedge clk); dir_r = 1; data_in = 75;
        @(posedge clk); dir_r = 1; data_in = 56;
        @(posedge clk); dir_r = 1; data_in = 69;
        @(posedge clk); dir_r = 0; data_in = 21;
        @(posedge clk); dir_r = 0; data_in = 579;
        @(posedge clk); dir_r = 0; data_in = 561;
        @(posedge clk); dir_r = 0; data_in = 839;
        @(posedge clk); dir_r = 0; data_in = 43;
        @(posedge clk); dir_r = 1; data_in = 43;
        @(posedge clk); dir_r = 1; data_in = 891;
        @(posedge clk); dir_r = 0; data_in = 91;
        @(posedge clk); dir_r = 1; data_in = 525;
        @(posedge clk); dir_r = 1; data_in = 26;
        @(posedge clk); dir_r = 1; data_in = 249;
        @(posedge clk); dir_r = 1; data_in = 66;
        @(posedge clk); dir_r = 0; data_in = 566;
        @(posedge clk); dir_r = 0; data_in = 10;
        @(posedge clk); dir_r = 1; data_in = 25;
        @(posedge clk); dir_r = 1; data_in = 93;
        @(posedge clk); dir_r = 0; data_in = 99;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 80;
        @(posedge clk); dir_r = 1; data_in = 80;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 1; data_in = 23;
        @(posedge clk); dir_r = 0; data_in = 58;
        @(posedge clk); dir_r = 0; data_in = 166;
        @(posedge clk); dir_r = 1; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 530;
        @(posedge clk); dir_r = 0; data_in = 64;
        @(posedge clk); dir_r = 0; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 1; data_in = 669;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 71;
        @(posedge clk); dir_r = 1; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 4;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 0; data_in = 545;
        @(posedge clk); dir_r = 0; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 81;
        @(posedge clk); dir_r = 0; data_in = 381;
        @(posedge clk); dir_r = 0; data_in = 51;
        @(posedge clk); dir_r = 1; data_in = 832;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 1; data_in = 982;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 34;
        @(posedge clk); dir_r = 1; data_in = 894;
        @(posedge clk); dir_r = 0; data_in = 90;
        @(posedge clk); dir_r = 1; data_in = 18;
        @(posedge clk); dir_r = 1; data_in = 93;
        @(posedge clk); dir_r = 0; data_in = 235;
        @(posedge clk); dir_r = 0; data_in = 97;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 0; data_in = 74;
        @(posedge clk); dir_r = 0; data_in = 658;
        @(posedge clk); dir_r = 1; data_in = 603;
        @(posedge clk); dir_r = 1; data_in = 29;
        @(posedge clk); dir_r = 0; data_in = 761;
        @(posedge clk); dir_r = 0; data_in = 168;
        @(posedge clk); dir_r = 0; data_in = 99;
        @(posedge clk); dir_r = 1; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 8;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 34;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 1; data_in = 36;
        @(posedge clk); dir_r = 1; data_in = 48;
        @(posedge clk); dir_r = 0; data_in = 12;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 0; data_in = 78;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 0; data_in = 65;
        @(posedge clk); dir_r = 0; data_in = 311;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 1; data_in = 89;
        @(posedge clk); dir_r = 0; data_in = 183;
        @(posedge clk); dir_r = 0; data_in = 96;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 64;
        @(posedge clk); dir_r = 1; data_in = 864;
        @(posedge clk); dir_r = 0; data_in = 15;
        @(posedge clk); dir_r = 0; data_in = 926;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 66;
        @(posedge clk); dir_r = 1; data_in = 81;
        @(posedge clk); dir_r = 0; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 397;
        @(posedge clk); dir_r = 0; data_in = 76;
        @(posedge clk); dir_r = 0; data_in = 36;
        @(posedge clk); dir_r = 1; data_in = 636;
        @(posedge clk); dir_r = 0; data_in = 596;
        @(posedge clk); dir_r = 1; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 96;
        @(posedge clk); dir_r = 1; data_in = 77;
        @(posedge clk); dir_r = 0; data_in = 74;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 76;
        @(posedge clk); dir_r = 1; data_in = 368;
        @(posedge clk); dir_r = 0; data_in = 798;
        @(posedge clk); dir_r = 0; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 51;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 0; data_in = 60;
        @(posedge clk); dir_r = 1; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 195;
        @(posedge clk); dir_r = 1; data_in = 54;
        @(posedge clk); dir_r = 0; data_in = 241;
        @(posedge clk); dir_r = 0; data_in = 311;
        @(posedge clk); dir_r = 0; data_in = 48;
        @(posedge clk); dir_r = 0; data_in = 976;
        @(posedge clk); dir_r = 0; data_in = 76;
        @(posedge clk); dir_r = 0; data_in = 12;
        @(posedge clk); dir_r = 0; data_in = 581;
        @(posedge clk); dir_r = 0; data_in = 907;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 0; data_in = 65;
        @(posedge clk); dir_r = 0; data_in = 58;
        @(posedge clk); dir_r = 0; data_in = 644;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 517;
        @(posedge clk); dir_r = 0; data_in = 308;
        @(posedge clk); dir_r = 1; data_in = 25;
        @(posedge clk); dir_r = 1; data_in = 59;
        @(posedge clk); dir_r = 0; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 43;
        @(posedge clk); dir_r = 1; data_in = 94;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 0; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 601;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 62;
        @(posedge clk); dir_r = 1; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 323;
        @(posedge clk); dir_r = 0; data_in = 6;
        @(posedge clk); dir_r = 0; data_in = 31;
        @(posedge clk); dir_r = 1; data_in = 58;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 918;
        @(posedge clk); dir_r = 1; data_in = 660;
        @(posedge clk); dir_r = 1; data_in = 86;
        @(posedge clk); dir_r = 0; data_in = 7;
        @(posedge clk); dir_r = 1; data_in = 35;
        @(posedge clk); dir_r = 1; data_in = 72;
        @(posedge clk); dir_r = 1; data_in = 32;
        @(posedge clk); dir_r = 0; data_in = 197;
        @(posedge clk); dir_r = 0; data_in = 35;
        @(posedge clk); dir_r = 0; data_in = 69;
        @(posedge clk); dir_r = 0; data_in = 32;
        @(posedge clk); dir_r = 0; data_in = 28;
        @(posedge clk); dir_r = 0; data_in = 71;
        @(posedge clk); dir_r = 0; data_in = 253;
        @(posedge clk); dir_r = 1; data_in = 78;
        @(posedge clk); dir_r = 1; data_in = 75;
        @(posedge clk); dir_r = 1; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 48;
        @(posedge clk); dir_r = 1; data_in = 43;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 1; data_in = 86;
        @(posedge clk); dir_r = 0; data_in = 286;
        @(posedge clk); dir_r = 1; data_in = 409;
        @(posedge clk); dir_r = 1; data_in = 91;
        @(posedge clk); dir_r = 1; data_in = 5;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 78;
        @(posedge clk); dir_r = 1; data_in = 33;
        @(posedge clk); dir_r = 1; data_in = 76;
        @(posedge clk); dir_r = 1; data_in = 91;
        @(posedge clk); dir_r = 1; data_in = 19;
        @(posedge clk); dir_r = 1; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 0; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 58;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 0; data_in = 17;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 0; data_in = 80;
        @(posedge clk); dir_r = 1; data_in = 33;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 1; data_in = 58;
        @(posedge clk); dir_r = 0; data_in = 456;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 1; data_in = 10;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 0; data_in = 31;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 30;
        @(posedge clk); dir_r = 1; data_in = 46;
        @(posedge clk); dir_r = 1; data_in = 354;
        @(posedge clk); dir_r = 1; data_in = 19;
        @(posedge clk); dir_r = 0; data_in = 89;
        @(posedge clk); dir_r = 0; data_in = 30;
        @(posedge clk); dir_r = 1; data_in = 91;
        @(posedge clk); dir_r = 0; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 577;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 1; data_in = 98;
        @(posedge clk); dir_r = 1; data_in = 5;
        @(posedge clk); dir_r = 1; data_in = 937;
        @(posedge clk); dir_r = 0; data_in = 60;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 76;
        @(posedge clk); dir_r = 0; data_in = 89;
        @(posedge clk); dir_r = 0; data_in = 89;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 0; data_in = 319;
        @(posedge clk); dir_r = 1; data_in = 26;
        @(posedge clk); dir_r = 1; data_in = 40;
        @(posedge clk); dir_r = 0; data_in = 14;
        @(posedge clk); dir_r = 0; data_in = 99;
        @(posedge clk); dir_r = 0; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 82;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 0; data_in = 3;
        @(posedge clk); dir_r = 1; data_in = 3;
        @(posedge clk); dir_r = 1; data_in = 844;
        @(posedge clk); dir_r = 1; data_in = 356;
        @(posedge clk); dir_r = 1; data_in = 10;
        @(posedge clk); dir_r = 0; data_in = 36;
        @(posedge clk); dir_r = 0; data_in = 74;
        @(posedge clk); dir_r = 1; data_in = 76;
        @(posedge clk); dir_r = 1; data_in = 37;
        @(posedge clk); dir_r = 0; data_in = 715;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 647;
        @(posedge clk); dir_r = 0; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 45;
        @(posedge clk); dir_r = 0; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 403;
        @(posedge clk); dir_r = 0; data_in = 17;
        @(posedge clk); dir_r = 0; data_in = 147;
        @(posedge clk); dir_r = 0; data_in = 24;
        @(posedge clk); dir_r = 1; data_in = 34;
        @(posedge clk); dir_r = 1; data_in = 37;
        @(posedge clk); dir_r = 1; data_in = 61;
        @(posedge clk); dir_r = 0; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 60;
        @(posedge clk); dir_r = 0; data_in = 40;
        @(posedge clk); dir_r = 0; data_in = 698;
        @(posedge clk); dir_r = 0; data_in = 946;
        @(posedge clk); dir_r = 1; data_in = 144;
        @(posedge clk); dir_r = 0; data_in = 48;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 78;
        @(posedge clk); dir_r = 0; data_in = 40;
        @(posedge clk); dir_r = 0; data_in = 49;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 80;
        @(posedge clk); dir_r = 0; data_in = 80;
        @(posedge clk); dir_r = 0; data_in = 180;
        @(posedge clk); dir_r = 0; data_in = 32;
        @(posedge clk); dir_r = 0; data_in = 12;
        @(posedge clk); dir_r = 1; data_in = 7;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 43;
        @(posedge clk); dir_r = 0; data_in = 43;
        @(posedge clk); dir_r = 1; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 99;
        @(posedge clk); dir_r = 0; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 0; data_in = 19;
        @(posedge clk); dir_r = 1; data_in = 36;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 0; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 56;
        @(posedge clk); dir_r = 0; data_in = 41;
        @(posedge clk); dir_r = 1; data_in = 30;
        @(posedge clk); dir_r = 0; data_in = 99;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 1; data_in = 30;
        @(posedge clk); dir_r = 0; data_in = 93;
        @(posedge clk); dir_r = 0; data_in = 39;
        @(posedge clk); dir_r = 1; data_in = 67;
        @(posedge clk); dir_r = 1; data_in = 80;
        @(posedge clk); dir_r = 1; data_in = 56;
        @(posedge clk); dir_r = 1; data_in = 723;
        @(posedge clk); dir_r = 1; data_in = 76;
        @(posedge clk); dir_r = 0; data_in = 60;
        @(posedge clk); dir_r = 0; data_in = 40;
        @(posedge clk); dir_r = 1; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 563;
        @(posedge clk); dir_r = 0; data_in = 37;
        @(posedge clk); dir_r = 0; data_in = 28;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 5;
        @(posedge clk); dir_r = 0; data_in = 46;
        @(posedge clk); dir_r = 0; data_in = 35;
        @(posedge clk); dir_r = 0; data_in = 11;
        @(posedge clk); dir_r = 1; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 27;
        @(posedge clk); dir_r = 1; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 13;
        @(posedge clk); dir_r = 1; data_in = 734;
        @(posedge clk); dir_r = 1; data_in = 85;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 1; data_in = 33;
        @(posedge clk); dir_r = 0; data_in = 74;
        @(posedge clk); dir_r = 0; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 414;
        @(posedge clk); dir_r = 1; data_in = 14;
        @(posedge clk); dir_r = 0; data_in = 91;
        @(posedge clk); dir_r = 0; data_in = 16;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 1;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 76;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 0; data_in = 33;
        @(posedge clk); dir_r = 1; data_in = 5;
        @(posedge clk); dir_r = 0; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 70;
        @(posedge clk); dir_r = 0; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 62;
        @(posedge clk); dir_r = 1; data_in = 38;
        @(posedge clk); dir_r = 0; data_in = 60;
        @(posedge clk); dir_r = 0; data_in = 40;
        @(posedge clk); dir_r = 0; data_in = 72;
        @(posedge clk); dir_r = 1; data_in = 72;
        @(posedge clk); dir_r = 1; data_in = 275;
        @(posedge clk); dir_r = 0; data_in = 4;
        @(posedge clk); dir_r = 0; data_in = 32;
        @(posedge clk); dir_r = 0; data_in = 572;
        @(posedge clk); dir_r = 1; data_in = 92;
        @(posedge clk); dir_r = 1; data_in = 38;
        @(posedge clk); dir_r = 1; data_in = 3;
        @(posedge clk); dir_r = 0; data_in = 86;
        @(posedge clk); dir_r = 0; data_in = 14;
        @(posedge clk); dir_r = 1; data_in = 36;
        @(posedge clk); dir_r = 1; data_in = 87;
        @(posedge clk); dir_r = 0; data_in = 165;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 0; data_in = 28;
        @(posedge clk); dir_r = 1; data_in = 85;
        @(posedge clk); dir_r = 1; data_in = 744;
        @(posedge clk); dir_r = 1; data_in = 199;
        @(posedge clk); dir_r = 0; data_in = 499;
        @(posedge clk); dir_r = 0; data_in = 320;
        @(posedge clk); dir_r = 0; data_in = 17;
        @(posedge clk); dir_r = 1; data_in = 383;
        @(posedge clk); dir_r = 0; data_in = 650;
        @(posedge clk); dir_r = 0; data_in = 1;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 1; data_in = 170;
        @(posedge clk); dir_r = 0; data_in = 82;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 1; data_in = 71;
        @(posedge clk); dir_r = 0; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 50;
        @(posedge clk); dir_r = 1; data_in = 40;
        @(posedge clk); dir_r = 1; data_in = 10;
        @(posedge clk); dir_r = 1; data_in = 74;
        @(posedge clk); dir_r = 1; data_in = 616;
        @(posedge clk); dir_r = 0; data_in = 56;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 0; data_in = 76;
        @(posedge clk); dir_r = 1; data_in = 676;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 929;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 56;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 0; data_in = 66;
        @(posedge clk); dir_r = 0; data_in = 76;
        @(posedge clk); dir_r = 0; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 649;
        @(posedge clk); dir_r = 1; data_in = 49;
        @(posedge clk); dir_r = 0; data_in = 619;
        @(posedge clk); dir_r = 0; data_in = 19;
        @(posedge clk); dir_r = 0; data_in = 52;
        @(posedge clk); dir_r = 1; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 85;
        @(posedge clk); dir_r = 0; data_in = 812;
        @(posedge clk); dir_r = 0; data_in = 730;
        @(posedge clk); dir_r = 0; data_in = 58;
        @(posedge clk); dir_r = 0; data_in = 72;
        @(posedge clk); dir_r = 1; data_in = 672;
        @(posedge clk); dir_r = 1; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 37;
        @(posedge clk); dir_r = 1; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 35;
        @(posedge clk); dir_r = 0; data_in = 135;
        @(posedge clk); dir_r = 1; data_in = 82;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 54;
        @(posedge clk); dir_r = 0; data_in = 43;
        @(posedge clk); dir_r = 0; data_in = 57;
        @(posedge clk); dir_r = 1; data_in = 18;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 0; data_in = 64;
        @(posedge clk); dir_r = 1; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 33;
        @(posedge clk); dir_r = 1; data_in = 76;
        @(posedge clk); dir_r = 1; data_in = 73;
        @(posedge clk); dir_r = 0; data_in = 333;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 4;
        @(posedge clk); dir_r = 0; data_in = 93;
        @(posedge clk); dir_r = 1; data_in = 369;
        @(posedge clk); dir_r = 0; data_in = 76;
        @(posedge clk); dir_r = 1; data_in = 34;
        @(posedge clk); dir_r = 0; data_in = 12;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 0; data_in = 195;
        @(posedge clk); dir_r = 0; data_in = 39;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 1; data_in = 723;
        @(posedge clk); dir_r = 0; data_in = 66;
        @(posedge clk); dir_r = 1; data_in = 743;
        @(posedge clk); dir_r = 0; data_in = 430;
        @(posedge clk); dir_r = 1; data_in = 55;
        @(posedge clk); dir_r = 0; data_in = 975;
        @(posedge clk); dir_r = 1; data_in = 50;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 0; data_in = 62;
        @(posedge clk); dir_r = 0; data_in = 43;
        @(posedge clk); dir_r = 1; data_in = 635;
        @(posedge clk); dir_r = 0; data_in = 2;
        @(posedge clk); dir_r = 0; data_in = 464;
        @(posedge clk); dir_r = 0; data_in = 64;
        @(posedge clk); dir_r = 1; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 746;
        @(posedge clk); dir_r = 0; data_in = 641;
        @(posedge clk); dir_r = 1; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 80;
        @(posedge clk); dir_r = 0; data_in = 209;
        @(posedge clk); dir_r = 1; data_in = 40;
        @(posedge clk); dir_r = 1; data_in = 722;
        @(posedge clk); dir_r = 0; data_in = 26;
        @(posedge clk); dir_r = 0; data_in = 8;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 8;
        @(posedge clk); dir_r = 1; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 0; data_in = 17;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 86;
        @(posedge clk); dir_r = 1; data_in = 517;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 51;
        @(posedge clk); dir_r = 1; data_in = 18;
        @(posedge clk); dir_r = 1; data_in = 10;
        @(posedge clk); dir_r = 1; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 77;
        @(posedge clk); dir_r = 0; data_in = 673;
        @(posedge clk); dir_r = 1; data_in = 5;
        @(posedge clk); dir_r = 1; data_in = 23;
        @(posedge clk); dir_r = 0; data_in = 99;
        @(posedge clk); dir_r = 1; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 83;
        @(posedge clk); dir_r = 0; data_in = 142;
        @(posedge clk); dir_r = 1; data_in = 51;
        @(posedge clk); dir_r = 0; data_in = 7;
        @(posedge clk); dir_r = 1; data_in = 69;
        @(posedge clk); dir_r = 0; data_in = 7;
        @(posedge clk); dir_r = 0; data_in = 77;
        @(posedge clk); dir_r = 0; data_in = 54;
        @(posedge clk); dir_r = 1; data_in = 72;
        @(posedge clk); dir_r = 1; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 0; data_in = 993;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 96;
        @(posedge clk); dir_r = 0; data_in = 41;
        @(posedge clk); dir_r = 0; data_in = 21;
        @(posedge clk); dir_r = 0; data_in = 85;
        @(posedge clk); dir_r = 0; data_in = 85;
        @(posedge clk); dir_r = 0; data_in = 65;
        @(posedge clk); dir_r = 0; data_in = 35;
        @(posedge clk); dir_r = 0; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 27;
        @(posedge clk); dir_r = 0; data_in = 46;
        @(posedge clk); dir_r = 0; data_in = 13;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 1; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 54;
        @(posedge clk); dir_r = 0; data_in = 69;
        @(posedge clk); dir_r = 0; data_in = 912;
        @(posedge clk); dir_r = 0; data_in = 15;
        @(posedge clk); dir_r = 0; data_in = 55;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 838;
        @(posedge clk); dir_r = 1; data_in = 34;
        @(posedge clk); dir_r = 1; data_in = 240;
        @(posedge clk); dir_r = 0; data_in = 41;
        @(posedge clk); dir_r = 1; data_in = 41;
        @(posedge clk); dir_r = 0; data_in = 95;
        @(posedge clk); dir_r = 1; data_in = 195;
        @(posedge clk); dir_r = 0; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 689;
        @(posedge clk); dir_r = 0; data_in = 510;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 0; data_in = 94;
        @(posedge clk); dir_r = 1; data_in = 73;
        @(posedge clk); dir_r = 0; data_in = 76;
        @(posedge clk); dir_r = 0; data_in = 24;
        @(posedge clk); dir_r = 0; data_in = 62;
        @(posedge clk); dir_r = 1; data_in = 62;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 412;
        @(posedge clk); dir_r = 1; data_in = 18;
        @(posedge clk); dir_r = 1; data_in = 45;
        @(posedge clk); dir_r = 0; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 80;
        @(posedge clk); dir_r = 1; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 50;
        @(posedge clk); dir_r = 1; data_in = 54;
        @(posedge clk); dir_r = 1; data_in = 56;
        @(posedge clk); dir_r = 1; data_in = 40;
        @(posedge clk); dir_r = 0; data_in = 22;
        @(posedge clk); dir_r = 1; data_in = 22;
        @(posedge clk); dir_r = 0; data_in = 35;
        @(posedge clk); dir_r = 0; data_in = 425;
        @(posedge clk); dir_r = 0; data_in = 96;
        @(posedge clk); dir_r = 1; data_in = 98;
        @(posedge clk); dir_r = 1; data_in = 78;
        @(posedge clk); dir_r = 1; data_in = 80;
        @(posedge clk); dir_r = 1; data_in = 420;
        @(posedge clk); dir_r = 0; data_in = 91;
        @(posedge clk); dir_r = 1; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 2;
        @(posedge clk); dir_r = 0; data_in = 17;
        @(posedge clk); dir_r = 0; data_in = 389;
        @(posedge clk); dir_r = 1; data_in = 206;
        @(posedge clk); dir_r = 0; data_in = 962;
        @(posedge clk); dir_r = 0; data_in = 71;
        @(posedge clk); dir_r = 1; data_in = 67;
        @(posedge clk); dir_r = 1; data_in = 666;
        @(posedge clk); dir_r = 1; data_in = 67;
        @(posedge clk); dir_r = 1; data_in = 362;
        @(posedge clk); dir_r = 1; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 90;
        @(posedge clk); dir_r = 1; data_in = 541;
        @(posedge clk); dir_r = 0; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 939;
        @(posedge clk); dir_r = 1; data_in = 62;
        @(posedge clk); dir_r = 0; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 7;
        @(posedge clk); dir_r = 0; data_in = 17;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 1; data_in = 85;
        @(posedge clk); dir_r = 0; data_in = 48;
        @(posedge clk); dir_r = 0; data_in = 3;
        @(posedge clk); dir_r = 0; data_in = 197;
        @(posedge clk); dir_r = 1; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 376;
        @(posedge clk); dir_r = 0; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 497;
        @(posedge clk); dir_r = 0; data_in = 733;
        @(posedge clk); dir_r = 0; data_in = 42;
        @(posedge clk); dir_r = 0; data_in = 839;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 1; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 5;
        @(posedge clk); dir_r = 1; data_in = 30;
        @(posedge clk); dir_r = 1; data_in = 456;
        @(posedge clk); dir_r = 1; data_in = 123;
        @(posedge clk); dir_r = 0; data_in = 52;
        @(posedge clk); dir_r = 1; data_in = 33;
        @(posedge clk); dir_r = 0; data_in = 85;
        @(posedge clk); dir_r = 1; data_in = 81;
        @(posedge clk); dir_r = 0; data_in = 46;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 1; data_in = 829;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 27;
        @(posedge clk); dir_r = 1; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 993;
        @(posedge clk); dir_r = 0; data_in = 57;
        @(posedge clk); dir_r = 0; data_in = 498;
        @(posedge clk); dir_r = 0; data_in = 77;
        @(posedge clk); dir_r = 1; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 1; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 60;
        @(posedge clk); dir_r = 1; data_in = 60;
        @(posedge clk); dir_r = 0; data_in = 18;
        @(posedge clk); dir_r = 1; data_in = 8;
        @(posedge clk); dir_r = 1; data_in = 75;
        @(posedge clk); dir_r = 1; data_in = 35;
        @(posedge clk); dir_r = 0; data_in = 32;
        @(posedge clk); dir_r = 1; data_in = 85;
        @(posedge clk); dir_r = 0; data_in = 36;
        @(posedge clk); dir_r = 1; data_in = 777;
        @(posedge clk); dir_r = 0; data_in = 93;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 795;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 1; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 139;
        @(posedge clk); dir_r = 1; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 54;
        @(posedge clk); dir_r = 0; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 559;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 10;
        @(posedge clk); dir_r = 1; data_in = 2;
        @(posedge clk); dir_r = 0; data_in = 12;
        @(posedge clk); dir_r = 1; data_in = 45;
        @(posedge clk); dir_r = 0; data_in = 63;
        @(posedge clk); dir_r = 1; data_in = 43;
        @(posedge clk); dir_r = 1; data_in = 475;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 0; data_in = 64;
        @(posedge clk); dir_r = 0; data_in = 33;
        @(posedge clk); dir_r = 0; data_in = 5;
        @(posedge clk); dir_r = 1; data_in = 5;
        @(posedge clk); dir_r = 0; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 51;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 0; data_in = 7;
        @(posedge clk); dir_r = 0; data_in = 60;
        @(posedge clk); dir_r = 1; data_in = 35;
        @(posedge clk); dir_r = 0; data_in = 54;
        @(posedge clk); dir_r = 1; data_in = 51;
        @(posedge clk); dir_r = 1; data_in = 72;
        @(posedge clk); dir_r = 0; data_in = 45;
        @(posedge clk); dir_r = 0; data_in = 19;
        @(posedge clk); dir_r = 1; data_in = 239;
        @(posedge clk); dir_r = 1; data_in = 61;
        @(posedge clk); dir_r = 1; data_in = 96;
        @(posedge clk); dir_r = 1; data_in = 67;
        @(posedge clk); dir_r = 0; data_in = 63;
        @(posedge clk); dir_r = 1; data_in = 78;
        @(posedge clk); dir_r = 1; data_in = 555;
        @(posedge clk); dir_r = 1; data_in = 54;
        @(posedge clk); dir_r = 1; data_in = 92;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 26;
        @(posedge clk); dir_r = 0; data_in = 64;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 94;
        @(posedge clk); dir_r = 0; data_in = 26;
        @(posedge clk); dir_r = 0; data_in = 74;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 23;
        @(posedge clk); dir_r = 1; data_in = 507;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 1; data_in = 8;
        @(posedge clk); dir_r = 1; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 93;
        @(posedge clk); dir_r = 1; data_in = 215;
        @(posedge clk); dir_r = 1; data_in = 50;
        @(posedge clk); dir_r = 0; data_in = 66;
        @(posedge clk); dir_r = 1; data_in = 666;
        @(posedge clk); dir_r = 1; data_in = 55;
        @(posedge clk); dir_r = 0; data_in = 81;
        @(posedge clk); dir_r = 0; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 68;
        @(posedge clk); dir_r = 0; data_in = 62;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 1; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 0; data_in = 65;
        @(posedge clk); dir_r = 1; data_in = 74;
        @(posedge clk); dir_r = 1; data_in = 986;
        @(posedge clk); dir_r = 0; data_in = 77;
        @(posedge clk); dir_r = 0; data_in = 423;
        @(posedge clk); dir_r = 0; data_in = 82;
        @(posedge clk); dir_r = 0; data_in = 10;
        @(posedge clk); dir_r = 1; data_in = 623;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 1; data_in = 94;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 692;
        @(posedge clk); dir_r = 1; data_in = 8;
        @(posedge clk); dir_r = 0; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 81;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 0; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 85;
        @(posedge clk); dir_r = 0; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 96;
        @(posedge clk); dir_r = 1; data_in = 93;
        @(posedge clk); dir_r = 0; data_in = 226;
        @(posedge clk); dir_r = 0; data_in = 860;
        @(posedge clk); dir_r = 0; data_in = 77;
        @(posedge clk); dir_r = 1; data_in = 50;
        @(posedge clk); dir_r = 0; data_in = 70;
        @(posedge clk); dir_r = 0; data_in = 45;
        @(posedge clk); dir_r = 0; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 22;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 0; data_in = 22;
        @(posedge clk); dir_r = 0; data_in = 371;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 34;
        @(posedge clk); dir_r = 0; data_in = 781;
        @(posedge clk); dir_r = 1; data_in = 3;
        @(posedge clk); dir_r = 1; data_in = 50;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 77;
        @(posedge clk); dir_r = 0; data_in = 16;
        @(posedge clk); dir_r = 1; data_in = 50;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 0; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 910;
        @(posedge clk); dir_r = 1; data_in = 282;
        @(posedge clk); dir_r = 1; data_in = 794;
        @(posedge clk); dir_r = 0; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 0; data_in = 970;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 99;
        @(posedge clk); dir_r = 1; data_in = 69;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 0; data_in = 41;
        @(posedge clk); dir_r = 1; data_in = 198;
        @(posedge clk); dir_r = 0; data_in = 24;
        @(posedge clk); dir_r = 1; data_in = 767;
        @(posedge clk); dir_r = 1; data_in = 3;
        @(posedge clk); dir_r = 1; data_in = 82;
        @(posedge clk); dir_r = 1; data_in = 30;
        @(posedge clk); dir_r = 1; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 1; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 96;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 1; data_in = 932;
        @(posedge clk); dir_r = 0; data_in = 77;
        @(posedge clk); dir_r = 0; data_in = 36;
        @(posedge clk); dir_r = 0; data_in = 113;
        @(posedge clk); dir_r = 1; data_in = 17;
        @(posedge clk); dir_r = 1; data_in = 912;
        @(posedge clk); dir_r = 0; data_in = 203;
        @(posedge clk); dir_r = 1; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 199;
        @(posedge clk); dir_r = 0; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 174;
        @(posedge clk); dir_r = 0; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 60;
        @(posedge clk); dir_r = 0; data_in = 32;
        @(posedge clk); dir_r = 1; data_in = 71;
        @(posedge clk); dir_r = 0; data_in = 17;
        @(posedge clk); dir_r = 0; data_in = 82;
        @(posedge clk); dir_r = 1; data_in = 19;
        @(posedge clk); dir_r = 0; data_in = 19;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 0; data_in = 16;
        @(posedge clk); dir_r = 0; data_in = 270;
        @(posedge clk); dir_r = 0; data_in = 97;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 88;
        @(posedge clk); dir_r = 0; data_in = 84;
        @(posedge clk); dir_r = 0; data_in = 16;
        @(posedge clk); dir_r = 0; data_in = 96;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 0; data_in = 94;
        @(posedge clk); dir_r = 1; data_in = 451;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 1; data_in = 22;
        @(posedge clk); dir_r = 0; data_in = 89;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 1; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 92;
        @(posedge clk); dir_r = 1; data_in = 8;
        @(posedge clk); dir_r = 0; data_in = 939;
        @(posedge clk); dir_r = 0; data_in = 33;
        @(posedge clk); dir_r = 1; data_in = 72;
        @(posedge clk); dir_r = 1; data_in = 38;
        @(posedge clk); dir_r = 1; data_in = 62;
        @(posedge clk); dir_r = 0; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 970;
        @(posedge clk); dir_r = 0; data_in = 3;
        @(posedge clk); dir_r = 0; data_in = 792;
        @(posedge clk); dir_r = 0; data_in = 94;
        @(posedge clk); dir_r = 1; data_in = 38;
        @(posedge clk); dir_r = 1; data_in = 56;
        @(posedge clk); dir_r = 0; data_in = 62;
        @(posedge clk); dir_r = 0; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 71;
        @(posedge clk); dir_r = 0; data_in = 40;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 1; data_in = 2;
        @(posedge clk); dir_r = 1; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 71;
        @(posedge clk); dir_r = 0; data_in = 668;
        @(posedge clk); dir_r = 0; data_in = 34;
        @(posedge clk); dir_r = 0; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 72;
        @(posedge clk); dir_r = 0; data_in = 62;
        @(posedge clk); dir_r = 0; data_in = 630;
        @(posedge clk); dir_r = 0; data_in = 52;
        @(posedge clk); dir_r = 1; data_in = 56;
        @(posedge clk); dir_r = 1; data_in = 813;
        @(posedge clk); dir_r = 0; data_in = 13;
        @(posedge clk); dir_r = 0; data_in = 3;
        @(posedge clk); dir_r = 1; data_in = 39;
        @(posedge clk); dir_r = 1; data_in = 81;
        @(posedge clk); dir_r = 0; data_in = 52;
        @(posedge clk); dir_r = 1; data_in = 433;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 0; data_in = 39;
        @(posedge clk); dir_r = 1; data_in = 220;
        @(posedge clk); dir_r = 1; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 93;
        @(posedge clk); dir_r = 1; data_in = 722;
        @(posedge clk); dir_r = 1; data_in = 78;
        @(posedge clk); dir_r = 1; data_in = 733;
        @(posedge clk); dir_r = 0; data_in = 36;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 1; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 575;
        @(posedge clk); dir_r = 1; data_in = 2;
        @(posedge clk); dir_r = 0; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 18;
        @(posedge clk); dir_r = 0; data_in = 91;
        @(posedge clk); dir_r = 1; data_in = 39;
        @(posedge clk); dir_r = 0; data_in = 577;
        @(posedge clk); dir_r = 1; data_in = 980;
        @(posedge clk); dir_r = 1; data_in = 932;
        @(posedge clk); dir_r = 0; data_in = 32;
        @(posedge clk); dir_r = 1; data_in = 634;
        @(posedge clk); dir_r = 1; data_in = 407;
        @(posedge clk); dir_r = 1; data_in = 201;
        @(posedge clk); dir_r = 1; data_in = 563;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 581;
        @(posedge clk); dir_r = 1; data_in = 5;
        @(posedge clk); dir_r = 0; data_in = 52;
        @(posedge clk); dir_r = 0; data_in = 42;
        @(posedge clk); dir_r = 0; data_in = 260;
        @(posedge clk); dir_r = 0; data_in = 819;
        @(posedge clk); dir_r = 0; data_in = 34;
        @(posedge clk); dir_r = 1; data_in = 613;
        @(posedge clk); dir_r = 1; data_in = 61;
        @(posedge clk); dir_r = 0; data_in = 12;
        @(posedge clk); dir_r = 0; data_in = 442;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 1;
        @(posedge clk); dir_r = 0; data_in = 25;
        @(posedge clk); dir_r = 1; data_in = 91;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 805;
        @(posedge clk); dir_r = 1; data_in = 151;
        @(posedge clk); dir_r = 0; data_in = 630;
        @(posedge clk); dir_r = 0; data_in = 3;
        @(posedge clk); dir_r = 1; data_in = 60;
        @(posedge clk); dir_r = 1; data_in = 690;
        @(posedge clk); dir_r = 1; data_in = 37;
        @(posedge clk); dir_r = 1; data_in = 54;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 95;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 1; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 13;
        @(posedge clk); dir_r = 0; data_in = 33;
        @(posedge clk); dir_r = 1; data_in = 850;
        @(posedge clk); dir_r = 0; data_in = 30;
        @(posedge clk); dir_r = 1; data_in = 80;
        @(posedge clk); dir_r = 0; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 246;
        @(posedge clk); dir_r = 1; data_in = 93;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 1; data_in = 83;
        @(posedge clk); dir_r = 0; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 2;
        @(posedge clk); dir_r = 1; data_in = 803;
        @(posedge clk); dir_r = 1; data_in = 451;
        @(posedge clk); dir_r = 1; data_in = 46;
        @(posedge clk); dir_r = 1; data_in = 55;
        @(posedge clk); dir_r = 0; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 1; data_in = 62;
        @(posedge clk); dir_r = 0; data_in = 62;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 0; data_in = 50;
        @(posedge clk); dir_r = 0; data_in = 5;
        @(posedge clk); dir_r = 0; data_in = 341;
        @(posedge clk); dir_r = 0; data_in = 60;
        @(posedge clk); dir_r = 1; data_in = 14;
        @(posedge clk); dir_r = 0; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 58;
        @(posedge clk); dir_r = 1; data_in = 53;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 0; data_in = 658;
        @(posedge clk); dir_r = 0; data_in = 58;
        @(posedge clk); dir_r = 1; data_in = 81;
        @(posedge clk); dir_r = 0; data_in = 65;
        @(posedge clk); dir_r = 0; data_in = 15;
        @(posedge clk); dir_r = 0; data_in = 65;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 89;
        @(posedge clk); dir_r = 1; data_in = 503;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 13;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 89;
        @(posedge clk); dir_r = 1; data_in = 497;
        @(posedge clk); dir_r = 1; data_in = 5;
        @(posedge clk); dir_r = 0; data_in = 179;
        @(posedge clk); dir_r = 1; data_in = 28;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 1; data_in = 25;
        @(posedge clk); dir_r = 1; data_in = 32;
        @(posedge clk); dir_r = 0; data_in = 33;
        @(posedge clk); dir_r = 0; data_in = 99;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 30;
        @(posedge clk); dir_r = 0; data_in = 278;
        @(posedge clk); dir_r = 1; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 97;
        @(posedge clk); dir_r = 1; data_in = 48;
        @(posedge clk); dir_r = 0; data_in = 48;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 0; data_in = 588;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 0; data_in = 34;
        @(posedge clk); dir_r = 0; data_in = 72;
        @(posedge clk); dir_r = 1; data_in = 13;
        @(posedge clk); dir_r = 1; data_in = 63;
        @(posedge clk); dir_r = 1; data_in = 189;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 1; data_in = 8;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 860;
        @(posedge clk); dir_r = 0; data_in = 445;
        @(posedge clk); dir_r = 0; data_in = 182;
        @(posedge clk); dir_r = 1; data_in = 68;
        @(posedge clk); dir_r = 0; data_in = 132;
        @(posedge clk); dir_r = 0; data_in = 51;
        @(posedge clk); dir_r = 0; data_in = 85;
        @(posedge clk); dir_r = 1; data_in = 2;
        @(posedge clk); dir_r = 0; data_in = 702;
        @(posedge clk); dir_r = 0; data_in = 30;
        @(posedge clk); dir_r = 0; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 190;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 0; data_in = 50;
        @(posedge clk); dir_r = 1; data_in = 599;
        @(posedge clk); dir_r = 0; data_in = 24;
        @(posedge clk); dir_r = 1; data_in = 58;
        @(posedge clk); dir_r = 1; data_in = 1;
        @(posedge clk); dir_r = 0; data_in = 18;
        @(posedge clk); dir_r = 0; data_in = 883;
        @(posedge clk); dir_r = 0; data_in = 384;
        @(posedge clk); dir_r = 0; data_in = 84;
        @(posedge clk); dir_r = 0; data_in = 72;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 1; data_in = 89;
        @(posedge clk); dir_r = 0; data_in = 84;
        @(posedge clk); dir_r = 0; data_in = 4;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 1; data_in = 777;
        @(posedge clk); dir_r = 1; data_in = 30;
        @(posedge clk); dir_r = 1; data_in = 2;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 1; data_in = 10;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 1; data_in = 622;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 0; data_in = 37;
        @(posedge clk); dir_r = 0; data_in = 50;
        @(posedge clk); dir_r = 1; data_in = 50;
        @(posedge clk); dir_r = 1; data_in = 3;
        @(posedge clk); dir_r = 0; data_in = 684;
        @(posedge clk); dir_r = 1; data_in = 60;
        @(posedge clk); dir_r = 1; data_in = 71;
        @(posedge clk); dir_r = 1; data_in = 50;
        @(posedge clk); dir_r = 1; data_in = 49;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 1; data_in = 8;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 49;
        @(posedge clk); dir_r = 1; data_in = 862;
        @(posedge clk); dir_r = 1; data_in = 73;
        @(posedge clk); dir_r = 0; data_in = 86;
        @(posedge clk); dir_r = 1; data_in = 308;
        @(posedge clk); dir_r = 0; data_in = 42;
        @(posedge clk); dir_r = 0; data_in = 666;
        @(posedge clk); dir_r = 1; data_in = 14;
        @(posedge clk); dir_r = 0; data_in = 96;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 17;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 0; data_in = 82;
        @(posedge clk); dir_r = 1; data_in = 82;
        @(posedge clk); dir_r = 1; data_in = 77;
        @(posedge clk); dir_r = 1; data_in = 223;
        @(posedge clk); dir_r = 1; data_in = 7;
        @(posedge clk); dir_r = 1; data_in = 18;
        @(posedge clk); dir_r = 0; data_in = 25;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 0; data_in = 67;
        @(posedge clk); dir_r = 0; data_in = 810;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 0; data_in = 96;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 165;
        @(posedge clk); dir_r = 0; data_in = 897;
        @(posedge clk); dir_r = 1; data_in = 91;
        @(posedge clk); dir_r = 1; data_in = 17;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 246;
        @(posedge clk); dir_r = 1; data_in = 540;
        @(posedge clk); dir_r = 1; data_in = 22;
        @(posedge clk); dir_r = 1; data_in = 64;
        @(posedge clk); dir_r = 0; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 0; data_in = 816;
        @(posedge clk); dir_r = 1; data_in = 5;
        @(posedge clk); dir_r = 1; data_in = 525;
        @(posedge clk); dir_r = 1; data_in = 56;
        @(posedge clk); dir_r = 1; data_in = 51;
        @(posedge clk); dir_r = 1; data_in = 853;
        @(posedge clk); dir_r = 1; data_in = 10;
        @(posedge clk); dir_r = 0; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 0; data_in = 796;
        @(posedge clk); dir_r = 0; data_in = 422;
        @(posedge clk); dir_r = 0; data_in = 193;
        @(posedge clk); dir_r = 1; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 40;
        @(posedge clk); dir_r = 0; data_in = 48;
        @(posedge clk); dir_r = 1; data_in = 75;
        @(posedge clk); dir_r = 1; data_in = 444;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 27;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 0; data_in = 88;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 616;
        @(posedge clk); dir_r = 0; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 591;
        @(posedge clk); dir_r = 0; data_in = 90;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 0; data_in = 95;
        @(posedge clk); dir_r = 1; data_in = 88;
        @(posedge clk); dir_r = 1; data_in = 135;
        @(posedge clk); dir_r = 0; data_in = 35;
        @(posedge clk); dir_r = 1; data_in = 96;
        @(posedge clk); dir_r = 0; data_in = 16;
        @(posedge clk); dir_r = 1; data_in = 71;
        @(posedge clk); dir_r = 1; data_in = 2;
        @(posedge clk); dir_r = 1; data_in = 847;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 68;
        @(posedge clk); dir_r = 0; data_in = 65;
        @(posedge clk); dir_r = 1; data_in = 76;
        @(posedge clk); dir_r = 0; data_in = 90;
        @(posedge clk); dir_r = 0; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 46;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 0; data_in = 772;
        @(posedge clk); dir_r = 0; data_in = 38;
        @(posedge clk); dir_r = 0; data_in = 36;
        @(posedge clk); dir_r = 1; data_in = 62;
        @(posedge clk); dir_r = 1; data_in = 94;
        @(posedge clk); dir_r = 1; data_in = 54;
        @(posedge clk); dir_r = 1; data_in = 738;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 0; data_in = 703;
        @(posedge clk); dir_r = 1; data_in = 69;
        @(posedge clk); dir_r = 0; data_in = 60;
        @(posedge clk); dir_r = 1; data_in = 89;
        @(posedge clk); dir_r = 1; data_in = 19;
        @(posedge clk); dir_r = 1; data_in = 22;
        @(posedge clk); dir_r = 0; data_in = 774;
        @(posedge clk); dir_r = 1; data_in = 4;
        @(posedge clk); dir_r = 0; data_in = 577;
        @(posedge clk); dir_r = 0; data_in = 94;
        @(posedge clk); dir_r = 0; data_in = 452;
        @(posedge clk); dir_r = 1; data_in = 76;
        @(posedge clk); dir_r = 0; data_in = 51;
        @(posedge clk); dir_r = 0; data_in = 5;
        @(posedge clk); dir_r = 1; data_in = 85;
        @(posedge clk); dir_r = 1; data_in = 18;
        @(posedge clk); dir_r = 0; data_in = 843;
        @(posedge clk); dir_r = 0; data_in = 36;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 0; data_in = 86;
        @(posedge clk); dir_r = 0; data_in = 647;
        @(posedge clk); dir_r = 0; data_in = 64;
        @(posedge clk); dir_r = 1; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 75;
        @(posedge clk); dir_r = 1; data_in = 2;
        @(posedge clk); dir_r = 0; data_in = 40;
        @(posedge clk); dir_r = 1; data_in = 40;
        @(posedge clk); dir_r = 0; data_in = 981;
        @(posedge clk); dir_r = 1; data_in = 8;
        @(posedge clk); dir_r = 0; data_in = 72;
        @(posedge clk); dir_r = 1; data_in = 80;
        @(posedge clk); dir_r = 0; data_in = 941;
        @(posedge clk); dir_r = 1; data_in = 3;
        @(posedge clk); dir_r = 1; data_in = 7;
        @(posedge clk); dir_r = 0; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 96;
        @(posedge clk); dir_r = 1; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 272;
        @(posedge clk); dir_r = 1; data_in = 52;
        @(posedge clk); dir_r = 0; data_in = 666;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 2;
        @(posedge clk); dir_r = 0; data_in = 2;
        @(posedge clk); dir_r = 1; data_in = 644;
        @(posedge clk); dir_r = 0; data_in = 49;
        @(posedge clk); dir_r = 0; data_in = 95;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 1; data_in = 36;
        @(posedge clk); dir_r = 1; data_in = 77;
        @(posedge clk); dir_r = 1; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 94;
        @(posedge clk); dir_r = 1; data_in = 96;
        @(posedge clk); dir_r = 0; data_in = 65;
        @(posedge clk); dir_r = 0; data_in = 31;
        @(posedge clk); dir_r = 0; data_in = 691;
        @(posedge clk); dir_r = 1; data_in = 91;
        @(posedge clk); dir_r = 1; data_in = 67;
        @(posedge clk); dir_r = 0; data_in = 67;
        @(posedge clk); dir_r = 1; data_in = 89;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 914;
        @(posedge clk); dir_r = 0; data_in = 681;
        @(posedge clk); dir_r = 1; data_in = 12;
        @(posedge clk); dir_r = 1; data_in = 95;
        @(posedge clk); dir_r = 1; data_in = 88;
        @(posedge clk); dir_r = 1; data_in = 56;
        @(posedge clk); dir_r = 1; data_in = 67;
        @(posedge clk); dir_r = 1; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 91;
        @(posedge clk); dir_r = 1; data_in = 89;
        @(posedge clk); dir_r = 0; data_in = 595;
        @(posedge clk); dir_r = 1; data_in = 56;
        @(posedge clk); dir_r = 1; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 64;
        @(posedge clk); dir_r = 1; data_in = 46;
        @(posedge clk); dir_r = 0; data_in = 74;
        @(posedge clk); dir_r = 0; data_in = 8;
        @(posedge clk); dir_r = 1; data_in = 92;
        @(posedge clk); dir_r = 1; data_in = 986;
        @(posedge clk); dir_r = 1; data_in = 128;
        @(posedge clk); dir_r = 1; data_in = 94;
        @(posedge clk); dir_r = 1; data_in = 13;
        @(posedge clk); dir_r = 0; data_in = 66;
        @(posedge clk); dir_r = 0; data_in = 38;
        @(posedge clk); dir_r = 1; data_in = 38;
        @(posedge clk); dir_r = 1; data_in = 53;
        @(posedge clk); dir_r = 1; data_in = 66;
        @(posedge clk); dir_r = 1; data_in = 34;
        @(posedge clk); dir_r = 0; data_in = 993;
        @(posedge clk); dir_r = 1; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 80;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 0; data_in = 82;
        @(posedge clk); dir_r = 1; data_in = 2;
        @(posedge clk); dir_r = 0; data_in = 3;
        @(posedge clk); dir_r = 1; data_in = 69;
        @(posedge clk); dir_r = 0; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 41;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 1; data_in = 88;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 0; data_in = 45;
        @(posedge clk); dir_r = 0; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 56;
        @(posedge clk); dir_r = 0; data_in = 54;
        @(posedge clk); dir_r = 1; data_in = 18;
        @(posedge clk); dir_r = 1; data_in = 61;
        @(posedge clk); dir_r = 0; data_in = 41;
        @(posedge clk); dir_r = 0; data_in = 775;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 0; data_in = 54;
        @(posedge clk); dir_r = 0; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 50;
        @(posedge clk); dir_r = 1; data_in = 78;
        @(posedge clk); dir_r = 1; data_in = 19;
        @(posedge clk); dir_r = 1; data_in = 54;
        @(posedge clk); dir_r = 0; data_in = 523;
        @(posedge clk); dir_r = 0; data_in = 31;
        @(posedge clk); dir_r = 0; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 0; data_in = 214;
        @(posedge clk); dir_r = 1; data_in = 40;
        @(posedge clk); dir_r = 0; data_in = 724;
        @(posedge clk); dir_r = 1; data_in = 634;
        @(posedge clk); dir_r = 0; data_in = 34;
        @(posedge clk); dir_r = 1; data_in = 99;
        @(posedge clk); dir_r = 1; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 50;
        @(posedge clk); dir_r = 0; data_in = 429;
        @(posedge clk); dir_r = 0; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 926;
        @(posedge clk); dir_r = 1; data_in = 74;
        @(posedge clk); dir_r = 1; data_in = 768;
        @(posedge clk); dir_r = 1; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 21;
        @(posedge clk); dir_r = 0; data_in = 77;
        @(posedge clk); dir_r = 0; data_in = 512;
        @(posedge clk); dir_r = 0; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 48;
        @(posedge clk); dir_r = 0; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 648;
        @(posedge clk); dir_r = 0; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 96;
        @(posedge clk); dir_r = 1; data_in = 503;
        @(posedge clk); dir_r = 0; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 677;
        @(posedge clk); dir_r = 0; data_in = 42;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 530;
        @(posedge clk); dir_r = 0; data_in = 685;
        @(posedge clk); dir_r = 1; data_in = 78;
        @(posedge clk); dir_r = 1; data_in = 60;
        @(posedge clk); dir_r = 0; data_in = 62;
        @(posedge clk); dir_r = 1; data_in = 379;
        @(posedge clk); dir_r = 0; data_in = 91;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 7;
        @(posedge clk); dir_r = 0; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 46;
        @(posedge clk); dir_r = 1; data_in = 183;
        @(posedge clk); dir_r = 1; data_in = 102;
        @(posedge clk); dir_r = 0; data_in = 25;
        @(posedge clk); dir_r = 0; data_in = 32;
        @(posedge clk); dir_r = 1; data_in = 57;
        @(posedge clk); dir_r = 1; data_in = 43;
        @(posedge clk); dir_r = 0; data_in = 26;
        @(posedge clk); dir_r = 1; data_in = 75;
        @(posedge clk); dir_r = 1; data_in = 50;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 288;
        @(posedge clk); dir_r = 0; data_in = 47;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 286;
        @(posedge clk); dir_r = 0; data_in = 486;
        @(posedge clk); dir_r = 1; data_in = 74;
        @(posedge clk); dir_r = 1; data_in = 626;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 90;
        @(posedge clk); dir_r = 0; data_in = 57;
        @(posedge clk); dir_r = 1; data_in = 58;
        @(posedge clk); dir_r = 0; data_in = 25;
        @(posedge clk); dir_r = 1; data_in = 10;
        @(posedge clk); dir_r = 0; data_in = 243;
        @(posedge clk); dir_r = 0; data_in = 51;
        @(posedge clk); dir_r = 1; data_in = 736;
        @(posedge clk); dir_r = 0; data_in = 51;
        @(posedge clk); dir_r = 0; data_in = 34;
        @(posedge clk); dir_r = 1; data_in = 5;
        @(posedge clk); dir_r = 1; data_in = 73;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 0; data_in = 38;
        @(posedge clk); dir_r = 0; data_in = 7;
        @(posedge clk); dir_r = 1; data_in = 92;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 1; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 1; data_in = 18;
        @(posedge clk); dir_r = 0; data_in = 584;
        @(posedge clk); dir_r = 0; data_in = 35;
        @(posedge clk); dir_r = 1; data_in = 77;
        @(posedge clk); dir_r = 0; data_in = 762;
        @(posedge clk); dir_r = 1; data_in = 62;
        @(posedge clk); dir_r = 0; data_in = 905;
        @(posedge clk); dir_r = 0; data_in = 76;
        @(posedge clk); dir_r = 0; data_in = 13;
        @(posedge clk); dir_r = 1; data_in = 294;
        @(posedge clk); dir_r = 1; data_in = 94;
        @(posedge clk); dir_r = 0; data_in = 49;
        @(posedge clk); dir_r = 0; data_in = 307;
        @(posedge clk); dir_r = 1; data_in = 62;
        @(posedge clk); dir_r = 1; data_in = 383;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 0; data_in = 67;
        @(posedge clk); dir_r = 0; data_in = 366;
        @(posedge clk); dir_r = 0; data_in = 184;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 58;
        @(posedge clk); dir_r = 0; data_in = 45;
        @(posedge clk); dir_r = 0; data_in = 54;
        @(posedge clk); dir_r = 1; data_in = 41;
        @(posedge clk); dir_r = 1; data_in = 161;
        @(posedge clk); dir_r = 1; data_in = 3;
        @(posedge clk); dir_r = 0; data_in = 64;
        @(posedge clk); dir_r = 0; data_in = 31;
        @(posedge clk); dir_r = 0; data_in = 17;
        @(posedge clk); dir_r = 1; data_in = 48;
        @(posedge clk); dir_r = 1; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 90;
        @(posedge clk); dir_r = 0; data_in = 63;
        @(posedge clk); dir_r = 1; data_in = 330;
        @(posedge clk); dir_r = 0; data_in = 51;
        @(posedge clk); dir_r = 1; data_in = 99;
        @(posedge clk); dir_r = 0; data_in = 78;
        @(posedge clk); dir_r = 1; data_in = 96;
        @(posedge clk); dir_r = 1; data_in = 33;
        @(posedge clk); dir_r = 0; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 60;
        @(posedge clk); dir_r = 0; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 976;
        @(posedge clk); dir_r = 1; data_in = 40;
        @(posedge clk); dir_r = 0; data_in = 99;
        @(posedge clk); dir_r = 0; data_in = 76;
        @(posedge clk); dir_r = 0; data_in = 34;
        @(posedge clk); dir_r = 1; data_in = 77;
        @(posedge clk); dir_r = 0; data_in = 68;
        @(posedge clk); dir_r = 0; data_in = 80;
        @(posedge clk); dir_r = 0; data_in = 433;
        @(posedge clk); dir_r = 1; data_in = 38;
        @(posedge clk); dir_r = 1; data_in = 34;
        @(posedge clk); dir_r = 0; data_in = 249;
        @(posedge clk); dir_r = 0; data_in = 85;
        @(posedge clk); dir_r = 0; data_in = 146;
        @(posedge clk); dir_r = 1; data_in = 8;
        @(posedge clk); dir_r = 1; data_in = 43;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 1; data_in = 14;
        @(posedge clk); dir_r = 1; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 62;
        @(posedge clk); dir_r = 0; data_in = 25;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 27;
        @(posedge clk); dir_r = 1; data_in = 462;
        @(posedge clk); dir_r = 1; data_in = 51;
        @(posedge clk); dir_r = 0; data_in = 43;
        @(posedge clk); dir_r = 0; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 956;
        @(posedge clk); dir_r = 1; data_in = 444;
        @(posedge clk); dir_r = 1; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 880;
        @(posedge clk); dir_r = 1; data_in = 25;
        @(posedge clk); dir_r = 1; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 57;
        @(posedge clk); dir_r = 1; data_in = 43;
        @(posedge clk); dir_r = 1; data_in = 30;
        @(posedge clk); dir_r = 0; data_in = 41;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 1; data_in = 8;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 0; data_in = 37;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 1; data_in = 133;
        @(posedge clk); dir_r = 0; data_in = 594;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 46;
        @(posedge clk); dir_r = 1; data_in = 135;
        @(posedge clk); dir_r = 0; data_in = 58;
        @(posedge clk); dir_r = 1; data_in = 55;
        @(posedge clk); dir_r = 0; data_in = 197;
        @(posedge clk); dir_r = 0; data_in = 614;
        @(posedge clk); dir_r = 0; data_in = 86;
        @(posedge clk); dir_r = 0; data_in = 5;
        @(posedge clk); dir_r = 1; data_in = 5;
        @(posedge clk); dir_r = 0; data_in = 2;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 15;
        @(posedge clk); dir_r = 0; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 83;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 17;
        @(posedge clk); dir_r = 0; data_in = 74;
        @(posedge clk); dir_r = 1; data_in = 986;
        @(posedge clk); dir_r = 1; data_in = 960;
        @(posedge clk); dir_r = 1; data_in = 45;
        @(posedge clk); dir_r = 0; data_in = 847;
        @(posedge clk); dir_r = 0; data_in = 870;
        @(posedge clk); dir_r = 1; data_in = 17;
        @(posedge clk); dir_r = 0; data_in = 71;
        @(posedge clk); dir_r = 1; data_in = 19;
        @(posedge clk); dir_r = 0; data_in = 56;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 1; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 1; data_in = 43;
        @(posedge clk); dir_r = 1; data_in = 88;
        @(posedge clk); dir_r = 0; data_in = 19;
        @(posedge clk); dir_r = 0; data_in = 36;
        @(posedge clk); dir_r = 0; data_in = 42;
        @(posedge clk); dir_r = 0; data_in = 25;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 66;
        @(posedge clk); dir_r = 0; data_in = 71;
        @(posedge clk); dir_r = 0; data_in = 763;
        @(posedge clk); dir_r = 0; data_in = 89;
        @(posedge clk); dir_r = 0; data_in = 8;
        @(posedge clk); dir_r = 0; data_in = 3;
        @(posedge clk); dir_r = 1; data_in = 13;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 0; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 36;
        @(posedge clk); dir_r = 1; data_in = 29;
        @(posedge clk); dir_r = 0; data_in = 49;
        @(posedge clk); dir_r = 0; data_in = 51;
        @(posedge clk); dir_r = 0; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 4;
        @(posedge clk); dir_r = 0; data_in = 96;
        @(posedge clk); dir_r = 1; data_in = 598;
        @(posedge clk); dir_r = 0; data_in = 534;
        @(posedge clk); dir_r = 1; data_in = 968;
        @(posedge clk); dir_r = 0; data_in = 784;
        @(posedge clk); dir_r = 0; data_in = 586;
        @(posedge clk); dir_r = 0; data_in = 71;
        @(posedge clk); dir_r = 1; data_in = 36;
        @(posedge clk); dir_r = 0; data_in = 94;
        @(posedge clk); dir_r = 0; data_in = 941;
        @(posedge clk); dir_r = 0; data_in = 77;
        @(posedge clk); dir_r = 1; data_in = 74;
        @(posedge clk); dir_r = 1; data_in = 143;
        @(posedge clk); dir_r = 0; data_in = 778;
        @(posedge clk); dir_r = 0; data_in = 58;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 56;
        @(posedge clk); dir_r = 1; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 86;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 1; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 72;
        @(posedge clk); dir_r = 1; data_in = 36;
        @(posedge clk); dir_r = 1; data_in = 546;
        @(posedge clk); dir_r = 1; data_in = 18;
        @(posedge clk); dir_r = 1; data_in = 25;
        @(posedge clk); dir_r = 0; data_in = 76;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 196;
        @(posedge clk); dir_r = 0; data_in = 30;
        @(posedge clk); dir_r = 1; data_in = 99;
        @(posedge clk); dir_r = 1; data_in = 25;
        @(posedge clk); dir_r = 0; data_in = 921;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 0; data_in = 215;
        @(posedge clk); dir_r = 0; data_in = 17;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 0; data_in = 34;
        @(posedge clk); dir_r = 0; data_in = 19;
        @(posedge clk); dir_r = 0; data_in = 56;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 0; data_in = 10;
        @(posedge clk); dir_r = 1; data_in = 22;
        @(posedge clk); dir_r = 0; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 34;
        @(posedge clk); dir_r = 0; data_in = 93;
        @(posedge clk); dir_r = 0; data_in = 48;
        @(posedge clk); dir_r = 0; data_in = 52;
        @(posedge clk); dir_r = 0; data_in = 76;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 62;
        @(posedge clk); dir_r = 1; data_in = 75;
        @(posedge clk); dir_r = 0; data_in = 437;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 25;
        @(posedge clk); dir_r = 0; data_in = 86;
        @(posedge clk); dir_r = 1; data_in = 52;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 84;
        @(posedge clk); dir_r = 0; data_in = 550;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 1; data_in = 346;
        @(posedge clk); dir_r = 1; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 7;
        @(posedge clk); dir_r = 1; data_in = 34;
        @(posedge clk); dir_r = 1; data_in = 120;
        @(posedge clk); dir_r = 1; data_in = 480;
        @(posedge clk); dir_r = 1; data_in = 223;
        @(posedge clk); dir_r = 0; data_in = 12;
        @(posedge clk); dir_r = 1; data_in = 51;
        @(posedge clk); dir_r = 1; data_in = 25;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 702;
        @(posedge clk); dir_r = 1; data_in = 99;
        @(posedge clk); dir_r = 0; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 87;
        @(posedge clk); dir_r = 0; data_in = 17;
        @(posedge clk); dir_r = 1; data_in = 46;
        @(posedge clk); dir_r = 0; data_in = 54;
        @(posedge clk); dir_r = 0; data_in = 88;
        @(posedge clk); dir_r = 0; data_in = 52;
        @(posedge clk); dir_r = 0; data_in = 48;
        @(posedge clk); dir_r = 0; data_in = 89;
        @(posedge clk); dir_r = 0; data_in = 430;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 99;
        @(posedge clk); dir_r = 1; data_in = 99;
        @(posedge clk); dir_r = 1; data_in = 40;
        @(posedge clk); dir_r = 1; data_in = 315;
        @(posedge clk); dir_r = 1; data_in = 45;
        @(posedge clk); dir_r = 0; data_in = 62;
        @(posedge clk); dir_r = 0; data_in = 38;
        @(posedge clk); dir_r = 1; data_in = 130;
        @(posedge clk); dir_r = 1; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 39;
        @(posedge clk); dir_r = 0; data_in = 88;
        @(posedge clk); dir_r = 0; data_in = 698;
        @(posedge clk); dir_r = 1; data_in = 62;
        @(posedge clk); dir_r = 0; data_in = 46;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 5;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 74;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 32;
        @(posedge clk); dir_r = 0; data_in = 67;
        @(posedge clk); dir_r = 0; data_in = 1;
        @(posedge clk); dir_r = 0; data_in = 759;
        @(posedge clk); dir_r = 0; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 181;
        @(posedge clk); dir_r = 0; data_in = 54;
        @(posedge clk); dir_r = 0; data_in = 96;
        @(posedge clk); dir_r = 1; data_in = 80;
        @(posedge clk); dir_r = 0; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 43;
        @(posedge clk); dir_r = 0; data_in = 74;
        @(posedge clk); dir_r = 1; data_in = 851;
        @(posedge clk); dir_r = 1; data_in = 49;
        @(posedge clk); dir_r = 0; data_in = 3;
        @(posedge clk); dir_r = 0; data_in = 29;
        @(posedge clk); dir_r = 0; data_in = 10;
        @(posedge clk); dir_r = 1; data_in = 22;
        @(posedge clk); dir_r = 0; data_in = 80;
        @(posedge clk); dir_r = 1; data_in = 69;
        @(posedge clk); dir_r = 0; data_in = 69;
        @(posedge clk); dir_r = 0; data_in = 17;
        @(posedge clk); dir_r = 1; data_in = 17;
        @(posedge clk); dir_r = 1; data_in = 709;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 1; data_in = 19;
        @(posedge clk); dir_r = 0; data_in = 19;
        @(posedge clk); dir_r = 1; data_in = 28;
        @(posedge clk); dir_r = 0; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 88;
        @(posedge clk); dir_r = 0; data_in = 55;
        @(posedge clk); dir_r = 0; data_in = 97;
        @(posedge clk); dir_r = 1; data_in = 3;
        @(posedge clk); dir_r = 1; data_in = 39;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 468;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 0; data_in = 8;
        @(posedge clk); dir_r = 1; data_in = 341;
        @(posedge clk); dir_r = 0; data_in = 69;
        @(posedge clk); dir_r = 1; data_in = 20;
        @(posedge clk); dir_r = 1; data_in = 64;
        @(posedge clk); dir_r = 0; data_in = 92;
        @(posedge clk); dir_r = 1; data_in = 23;
        @(posedge clk); dir_r = 0; data_in = 8;
        @(posedge clk); dir_r = 1; data_in = 69;
        @(posedge clk); dir_r = 0; data_in = 47;
        @(posedge clk); dir_r = 1; data_in = 64;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 71;
        @(posedge clk); dir_r = 1; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 1; data_in = 7;
        @(posedge clk); dir_r = 0; data_in = 7;
        @(posedge clk); dir_r = 0; data_in = 292;
        @(posedge clk); dir_r = 0; data_in = 93;
        @(posedge clk); dir_r = 1; data_in = 584;
        @(posedge clk); dir_r = 1; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 1; data_in = 94;
        @(posedge clk); dir_r = 0; data_in = 69;
        @(posedge clk); dir_r = 0; data_in = 15;
        @(posedge clk); dir_r = 0; data_in = 379;
        @(posedge clk); dir_r = 0; data_in = 6;
        @(posedge clk); dir_r = 0; data_in = 621;
        @(posedge clk); dir_r = 1; data_in = 3;
        @(posedge clk); dir_r = 0; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 97;
        @(posedge clk); dir_r = 1; data_in = 57;
        @(posedge clk); dir_r = 0; data_in = 357;
        @(posedge clk); dir_r = 0; data_in = 82;
        @(posedge clk); dir_r = 1; data_in = 533;
        @(posedge clk); dir_r = 0; data_in = 71;
        @(posedge clk); dir_r = 0; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 0; data_in = 84;
        @(posedge clk); dir_r = 0; data_in = 60;
        @(posedge clk); dir_r = 1; data_in = 598;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 1; data_in = 523;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 0; data_in = 780;
        @(posedge clk); dir_r = 0; data_in = 420;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 753;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 42;
        @(posedge clk); dir_r = 0; data_in = 78;
        @(posedge clk); dir_r = 0; data_in = 40;
        @(posedge clk); dir_r = 1; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 77;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 1; data_in = 682;
        @(posedge clk); dir_r = 0; data_in = 25;
        @(posedge clk); dir_r = 0; data_in = 875;
        @(posedge clk); dir_r = 1; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 32;
        @(posedge clk); dir_r = 0; data_in = 71;
        @(posedge clk); dir_r = 0; data_in = 43;
        @(posedge clk); dir_r = 1; data_in = 14;
        @(posedge clk); dir_r = 0; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 13;
        @(posedge clk); dir_r = 0; data_in = 89;
        @(posedge clk); dir_r = 1; data_in = 60;
        @(posedge clk); dir_r = 1; data_in = 22;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 83;
        @(posedge clk); dir_r = 0; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 63;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 0; data_in = 36;
        @(posedge clk); dir_r = 1; data_in = 95;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 403;
        @(posedge clk); dir_r = 1; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 14;
        @(posedge clk); dir_r = 0; data_in = 90;
        @(posedge clk); dir_r = 1; data_in = 251;
        @(posedge clk); dir_r = 0; data_in = 99;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 575;
        @(posedge clk); dir_r = 1; data_in = 66;
        @(posedge clk); dir_r = 1; data_in = 840;
        @(posedge clk); dir_r = 1; data_in = 23;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 1; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 39;
        @(posedge clk); dir_r = 0; data_in = 5;
        @(posedge clk); dir_r = 1; data_in = 614;
        @(posedge clk); dir_r = 1; data_in = 390;
        @(posedge clk); dir_r = 0; data_in = 22;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 1; data_in = 256;
        @(posedge clk); dir_r = 0; data_in = 889;
        @(posedge clk); dir_r = 1; data_in = 32;
        @(posedge clk); dir_r = 1; data_in = 57;
        @(posedge clk); dir_r = 0; data_in = 83;
        @(posedge clk); dir_r = 1; data_in = 7;
        @(posedge clk); dir_r = 1; data_in = 876;
        @(posedge clk); dir_r = 0; data_in = 10;
        @(posedge clk); dir_r = 1; data_in = 74;
        @(posedge clk); dir_r = 0; data_in = 74;
        @(posedge clk); dir_r = 0; data_in = 91;
        @(posedge clk); dir_r = 0; data_in = 57;
        @(posedge clk); dir_r = 0; data_in = 69;
        @(posedge clk); dir_r = 0; data_in = 40;
        @(posedge clk); dir_r = 0; data_in = 76;
        @(posedge clk); dir_r = 1; data_in = 86;
        @(posedge clk); dir_r = 1; data_in = 393;
        @(posedge clk); dir_r = 1; data_in = 64;
        @(posedge clk); dir_r = 1; data_in = 22;
        @(posedge clk); dir_r = 0; data_in = 22;
        @(posedge clk); dir_r = 1; data_in = 10;
        @(posedge clk); dir_r = 1; data_in = 13;
        @(posedge clk); dir_r = 1; data_in = 63;
        @(posedge clk); dir_r = 0; data_in = 80;
        @(posedge clk); dir_r = 0; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 195;
        @(posedge clk); dir_r = 1; data_in = 38;
        @(posedge clk); dir_r = 1; data_in = 67;
        @(posedge clk); dir_r = 0; data_in = 57;
        @(posedge clk); dir_r = 1; data_in = 26;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 0; data_in = 158;
        @(posedge clk); dir_r = 0; data_in = 883;
        @(posedge clk); dir_r = 1; data_in = 104;
        @(posedge clk); dir_r = 1; data_in = 37;
        @(posedge clk); dir_r = 0; data_in = 41;
        @(posedge clk); dir_r = 0; data_in = 5;
        @(posedge clk); dir_r = 1; data_in = 69;
        @(posedge clk); dir_r = 0; data_in = 970;
        @(posedge clk); dir_r = 0; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 245;
        @(posedge clk); dir_r = 1; data_in = 982;
        @(posedge clk); dir_r = 1; data_in = 418;
        @(posedge clk); dir_r = 1; data_in = 67;
        @(posedge clk); dir_r = 0; data_in = 67;
        @(posedge clk); dir_r = 1; data_in = 247;
        @(posedge clk); dir_r = 1; data_in = 19;
        @(posedge clk); dir_r = 1; data_in = 34;
        @(posedge clk); dir_r = 1; data_in = 934;
        @(posedge clk); dir_r = 0; data_in = 922;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 1; data_in = 59;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 0; data_in = 20;
        @(posedge clk); dir_r = 0; data_in = 80;
        @(posedge clk); dir_r = 0; data_in = 817;
        @(posedge clk); dir_r = 0; data_in = 10;
        @(posedge clk); dir_r = 0; data_in = 818;
        @(posedge clk); dir_r = 0; data_in = 55;
        @(posedge clk); dir_r = 0; data_in = 552;
        @(posedge clk); dir_r = 1; data_in = 87;
        @(posedge clk); dir_r = 1; data_in = 875;
        @(posedge clk); dir_r = 0; data_in = 10;
        @(posedge clk); dir_r = 0; data_in = 935;
        @(posedge clk); dir_r = 0; data_in = 18;
        @(posedge clk); dir_r = 0; data_in = 47;
        @(posedge clk); dir_r = 1; data_in = 50;
        @(posedge clk); dir_r = 0; data_in = 50;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 1; data_in = 91;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 1; data_in = 553;
        @(posedge clk); dir_r = 0; data_in = 29;
        @(posedge clk); dir_r = 0; data_in = 71;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 0; data_in = 11;
        @(posedge clk); dir_r = 1; data_in = 10;
        @(posedge clk); dir_r = 0; data_in = 90;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 322;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 51;
        @(posedge clk); dir_r = 1; data_in = 38;
        @(posedge clk); dir_r = 0; data_in = 115;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 0; data_in = 13;
        @(posedge clk); dir_r = 1; data_in = 72;
        @(posedge clk); dir_r = 1; data_in = 99;
        @(posedge clk); dir_r = 1; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 1; data_in = 58;
        @(posedge clk); dir_r = 1; data_in = 33;
        @(posedge clk); dir_r = 1; data_in = 384;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 1; data_in = 72;
        @(posedge clk); dir_r = 0; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 372;
        @(posedge clk); dir_r = 1; data_in = 51;
        @(posedge clk); dir_r = 0; data_in = 62;
        @(posedge clk); dir_r = 1; data_in = 21;
        @(posedge clk); dir_r = 0; data_in = 15;
        @(posedge clk); dir_r = 0; data_in = 743;
        @(posedge clk); dir_r = 0; data_in = 206;
        @(posedge clk); dir_r = 1; data_in = 64;
        @(posedge clk); dir_r = 0; data_in = 22;
        @(posedge clk); dir_r = 0; data_in = 90;
        @(posedge clk); dir_r = 0; data_in = 14;
        @(posedge clk); dir_r = 1; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 72;
        @(posedge clk); dir_r = 0; data_in = 55;
        @(posedge clk); dir_r = 1; data_in = 65;
        @(posedge clk); dir_r = 0; data_in = 10;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 0; data_in = 71;
        @(posedge clk); dir_r = 0; data_in = 26;
        @(posedge clk); dir_r = 1; data_in = 4;
        @(posedge clk); dir_r = 0; data_in = 66;
        @(posedge clk); dir_r = 0; data_in = 72;
        @(posedge clk); dir_r = 1; data_in = 46;
        @(posedge clk); dir_r = 1; data_in = 523;
        @(posedge clk); dir_r = 1; data_in = 751;
        @(posedge clk); dir_r = 0; data_in = 28;
        @(posedge clk); dir_r = 1; data_in = 560;
        @(posedge clk); dir_r = 0; data_in = 52;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 1; data_in = 81;
        @(posedge clk); dir_r = 0; data_in = 158;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 853;
        @(posedge clk); dir_r = 0; data_in = 820;
        @(posedge clk); dir_r = 0; data_in = 13;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 41;
        @(posedge clk); dir_r = 0; data_in = 292;
        @(posedge clk); dir_r = 0; data_in = 34;
        @(posedge clk); dir_r = 0; data_in = 827;
        @(posedge clk); dir_r = 0; data_in = 99;
        @(posedge clk); dir_r = 0; data_in = 937;
        @(posedge clk); dir_r = 0; data_in = 37;
        @(posedge clk); dir_r = 1; data_in = 94;
        @(posedge clk); dir_r = 0; data_in = 94;
        @(posedge clk); dir_r = 1; data_in = 73;
        @(posedge clk); dir_r = 0; data_in = 41;
        @(posedge clk); dir_r = 0; data_in = 607;
        @(posedge clk); dir_r = 0; data_in = 25;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 0; data_in = 6;
        @(posedge clk); dir_r = 0; data_in = 26;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 88;
        @(posedge clk); dir_r = 0; data_in = 56;
        @(posedge clk); dir_r = 0; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 27;
        @(posedge clk); dir_r = 1; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 10;
        @(posedge clk); dir_r = 0; data_in = 10;
        @(posedge clk); dir_r = 1; data_in = 94;
        @(posedge clk); dir_r = 0; data_in = 28;
        @(posedge clk); dir_r = 1; data_in = 46;
        @(posedge clk); dir_r = 0; data_in = 39;
        @(posedge clk); dir_r = 0; data_in = 402;
        @(posedge clk); dir_r = 1; data_in = 59;
        @(posedge clk); dir_r = 0; data_in = 425;
        @(posedge clk); dir_r = 1; data_in = 195;
        @(posedge clk); dir_r = 1; data_in = 51;
        @(posedge clk); dir_r = 0; data_in = 51;
        @(posedge clk); dir_r = 1; data_in = 58;
        @(posedge clk); dir_r = 0; data_in = 8;
        @(posedge clk); dir_r = 1; data_in = 50;
        @(posedge clk); dir_r = 0; data_in = 5;
        @(posedge clk); dir_r = 0; data_in = 404;
        @(posedge clk); dir_r = 0; data_in = 91;
        @(posedge clk); dir_r = 0; data_in = 14;
        @(posedge clk); dir_r = 1; data_in = 14;
        @(posedge clk); dir_r = 1; data_in = 56;
        @(posedge clk); dir_r = 0; data_in = 56;
        @(posedge clk); dir_r = 0; data_in = 33;
        @(posedge clk); dir_r = 0; data_in = 67;
        @(posedge clk); dir_r = 0; data_in = 98;
        @(posedge clk); dir_r = 0; data_in = 45;
        @(posedge clk); dir_r = 1; data_in = 85;
        @(posedge clk); dir_r = 0; data_in = 42;
        @(posedge clk); dir_r = 1; data_in = 41;
        @(posedge clk); dir_r = 1; data_in = 26;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 54;
        @(posedge clk); dir_r = 0; data_in = 225;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 0; data_in = 17;
        @(posedge clk); dir_r = 0; data_in = 22;
        @(posedge clk); dir_r = 1; data_in = 94;
        @(posedge clk); dir_r = 1; data_in = 10;
        @(posedge clk); dir_r = 1; data_in = 510;
        @(posedge clk); dir_r = 1; data_in = 80;
        @(posedge clk); dir_r = 0; data_in = 22;
        @(posedge clk); dir_r = 1; data_in = 60;
        @(posedge clk); dir_r = 0; data_in = 47;
        @(posedge clk); dir_r = 1; data_in = 36;
        @(posedge clk); dir_r = 0; data_in = 127;
        @(posedge clk); dir_r = 0; data_in = 163;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 0; data_in = 52;
        @(posedge clk); dir_r = 0; data_in = 96;
        @(posedge clk); dir_r = 1; data_in = 70;
        @(posedge clk); dir_r = 1; data_in = 53;
        @(posedge clk); dir_r = 1; data_in = 73;
        @(posedge clk); dir_r = 1; data_in = 91;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 33;
        @(posedge clk); dir_r = 1; data_in = 33;
        @(posedge clk); dir_r = 1; data_in = 14;
        @(posedge clk); dir_r = 1; data_in = 39;
        @(posedge clk); dir_r = 0; data_in = 53;
        @(posedge clk); dir_r = 1; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 76;
        @(posedge clk); dir_r = 1; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 1;
        @(posedge clk); dir_r = 1; data_in = 60;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 1; data_in = 51;
        @(posedge clk); dir_r = 1; data_in = 39;
        @(posedge clk); dir_r = 1; data_in = 68;
        @(posedge clk); dir_r = 1; data_in = 7;
        @(posedge clk); dir_r = 1; data_in = 29;
        @(posedge clk); dir_r = 0; data_in = 43;
        @(posedge clk); dir_r = 1; data_in = 88;
        @(posedge clk); dir_r = 0; data_in = 22;
        @(posedge clk); dir_r = 0; data_in = 31;
        @(posedge clk); dir_r = 0; data_in = 5;
        @(posedge clk); dir_r = 0; data_in = 30;
        @(posedge clk); dir_r = 0; data_in = 99;
        @(posedge clk); dir_r = 0; data_in = 84;
        @(posedge clk); dir_r = 1; data_in = 79;
        @(posedge clk); dir_r = 0; data_in = 72;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 30;
        @(posedge clk); dir_r = 0; data_in = 28;
        @(posedge clk); dir_r = 1; data_in = 59;
        @(posedge clk); dir_r = 1; data_in = 41;
        @(posedge clk); dir_r = 0; data_in = 82;
        @(posedge clk); dir_r = 0; data_in = 34;
        @(posedge clk); dir_r = 1; data_in = 34;
        @(posedge clk); dir_r = 0; data_in = 24;
        @(posedge clk); dir_r = 0; data_in = 79;
        @(posedge clk); dir_r = 1; data_in = 54;
        @(posedge clk); dir_r = 1; data_in = 49;
        @(posedge clk); dir_r = 1; data_in = 95;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 90;
        @(posedge clk); dir_r = 0; data_in = 61;
        @(posedge clk); dir_r = 0; data_in = 39;
        @(posedge clk); dir_r = 0; data_in = 14;
        @(posedge clk); dir_r = 1; data_in = 14;
        @(posedge clk); dir_r = 1; data_in = 8;
        @(posedge clk); dir_r = 1; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 34;
        @(posedge clk); dir_r = 1; data_in = 16;
        @(posedge clk); dir_r = 0; data_in = 14;
        @(posedge clk); dir_r = 1; data_in = 28;
        @(posedge clk); dir_r = 1; data_in = 46;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 1; data_in = 22;
        @(posedge clk); dir_r = 1; data_in = 30;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 0; data_in = 4;
        @(posedge clk); dir_r = 1; data_in = 35;
        @(posedge clk); dir_r = 1; data_in = 48;
        @(posedge clk); dir_r = 0; data_in = 39;
        @(posedge clk); dir_r = 0; data_in = 15;
        @(posedge clk); dir_r = 1; data_in = 46;
        @(posedge clk); dir_r = 1; data_in = 34;
        @(posedge clk); dir_r = 0; data_in = 11;
        @(posedge clk); dir_r = 1; data_in = 17;
        @(posedge clk); dir_r = 1; data_in = 10;
        @(posedge clk); dir_r = 1; data_in = 24;
        @(posedge clk); dir_r = 1; data_in = 31;
        @(posedge clk); dir_r = 1; data_in = 18;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 5;
        @(posedge clk); dir_r = 1; data_in = 38;
        @(posedge clk); dir_r = 0; data_in = 3;
        @(posedge clk); dir_r = 0; data_in = 27;
        @(posedge clk); dir_r = 0; data_in = 7;
        @(posedge clk); dir_r = 0; data_in = 30;
        @(posedge clk); dir_r = 0; data_in = 10;
        @(posedge clk); dir_r = 0; data_in = 2;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 6;
        @(posedge clk); dir_r = 1; data_in = 5;
        @(posedge clk); dir_r = 0; data_in = 46;
        @(posedge clk); dir_r = 1; data_in = 15;
        @(posedge clk); dir_r = 0; data_in = 44;
        @(posedge clk); dir_r = 1; data_in = 33;
        @(posedge clk); dir_r = 1; data_in = 11;
        @(posedge clk); dir_r = 0; data_in = 9;
        @(posedge clk); dir_r = 0; data_in = 23;
        @(posedge clk); dir_r = 1; data_in = 30;
        @(posedge clk); dir_r = 1; data_in = 29;
        @(posedge clk); dir_r = 1; data_in = 47;
        @(posedge clk); dir_r = 0; data_in = 34;
        // === END INPUT SEQUENCE ===

        // Print final result
        #20;
        $display("=== TEST COMPLETE ===");
        $display("Final zero_count = %d", zero_count);
        $display("Final zero_cros = %d", zero_cross);

        $finish;
    end

endmodule

