module hardware_wrapper(
    
)

endmodule